--------------------------------------------------------------------------------
-- Engineer:  Luca Caronti    [luca.caronti@studenti.unit.it]
--            Simone Ruffini  [simone.ruffini@tutanota.com]
--
-- Create Date:   05/17/2020 03:21:54 PM
-- Design Name:
-- Module Name:   INT_EMU - Behavioral
-- Project Name:  NORM
--
-- Description: Intermittency emulation core.
-- Details: This entity generates a signal (RST_EMU) used by the test platform
--  as a reset signal. This is generated by comparing a voltage sample to a
--  voltage level selected as the reset threshold.
--
-- Revision:
-- Revision 00 - Luca Caronti
-- * file created
-- Revision 01 - Simone Ruffini
-- * refactoring and generalizatin of the component (input rom is outside of the entity)
-- Additional Comments:
--
--------------------------------------------------------------------------------

----------------------------- PACKAGES/LIBRARIES -------------------------------

library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.NUMERIC_STD.all;

  -- User libraries
  use work.NORM_PKG.all;

----------------------------- ENTITY -------------------------------------------

entity INT_EMU is
  generic (
    VTRACE_ROM_NUM_ELEMENTS     : natural;                                                     -- Number of samples inside of Voltage Trace ROM
    NUM_THRESHOLDS              : natural := 1;                                                -- Number of compared thresholds (the one for RST_EMU is one too)
    SAMPLES_PRESCALER           : natural := 1                                                 -- Sampling from ROM prescaler value (NOTE: > 0)
  );
  port (
    CLK                         : in    std_logic;                                                -- Clock signal
    RST                         : in    std_logic;                                                -- Positive reset
    EN                          : in    std_logic;                                                -- Enable core
    INIT                        : in    std_logic;                                                -- Init core
    RST_EMU                     : out   std_logic;                                                -- Emulated positive reset
    THRESH_STATS                : out   std_logic_vector(NUM_THRESHOLDS - 1 downto 0);            -- Thresholds statuses
    THRESH_VALUES               : in    thresh_values_t(NUM_THRESHOLDS - 1 downto 0);             -- Thresholds values
    RST_EMU_THRESH_INDX         : in    natural range 0 to NUM_THRESHOLDS - 1;                    -- Index of threshold used for RST_EMU
    VTRACE_ROM_START_INDX       : in    natural;                                                  -- Voltage Trace ROM sampling start index
    VTRACE_ROM_SAMPLES          : in    natural;                                                  -- Voltage Trace ROM number of used samples from VTRACE_ROM_START_INDX
    VTRACE_ROM_RADDR            : out   natural;                                                  -- ROM read address
    VTRACE_ROM_DOUT             : in    integer                                                   -- ROM data output
  );
end entity INT_EMU;

----------------------------- ARCHITECTURE -------------------------------------

architecture BEHAVIORAL of INT_EMU is

  --########################### CONSTANTS 1 ####################################

  --########################### TYPES ##########################################

  --########################### FUNCTIONS ######################################

  --########################### CONSTANTS 2 ####################################

  --########################### SIGNALS ########################################

  signal rst_emu_s             : std_logic;
  signal rst_emu_gate          : std_logic := '0';
  signal rom_start_addr_samp   : natural := 0;
  signal rom_offset_samp       : natural := 0;
  signal rom_raddr_s           : natural := 0;
  signal output_comparator     : std_logic_vector(NUM_THRESHOLDS - 1 downto 0);
  signal prescaler_cnt_tc      : std_logic;
  signal prescaler_cnt_init    : std_logic;

  --########################### ARCHITECTURE BEGIN #############################

begin

  assert (SAMPLES_PRESCALER > 0)
    report "The prescaler for the sampling time must be greater then 0"
    severity failure;

  --########################### ENTITY DEFINITION ##############################

  U_PRESCALER : entity work.cnt
    generic map (
      MAX         => SAMPLES_PRESCALER - 1,
      INIT_VALUE  => SAMPLES_PRESCALER - 1,
      INCREASE_BY => 1
    )
    port map (
      CLK   => CLK,
      RST   => RST,
      INIT  => prescaler_cnt_init,
      CE    => '1',
      TC    => prescaler_cnt_tc,
      VALUE => open
    );

  --########################## OUTPUT PORTS WIRING #############################

  RST_EMU <= rst_emu_s;

  THRESH_STATS <= output_comparator;

  VTRACE_ROM_RADDR <= rom_raddr_s;

  --########################## COBINATORIAL FUNCTIONS ##########################

  G_COMPARATOR : for i in NUM_THRESHOLDS - 1  downto 0 generate
    output_comparator(i) <= '1' when VTRACE_ROM_DOUT <= THRESH_VALUES(i) else
                            '0';
  end generate G_COMPARATOR;

  rst_emu_s <= (rst_emu_gate AND output_comparator(RST_EMU_THRESH_INDX)) OR RST;

  --########################## PROCESSES #######################################

  --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
  -- Init Delay
  --
  -- Keep init signal after rst is down for the rest of the clock cycle
  -- this lets PRESCALER_CNT more init time

  P_INIT_DELAY : process (CLK) is
  begin

    if (CLK'event and CLK = '1') then
      prescaler_cnt_init <= '0';
      if (RST = '1') then
        prescaler_cnt_init <= '1';
      end if;
    end if;

  end process P_INIT_DELAY;

  --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
  -- Samples rom start address and rom offset
  --
  -- These signals can change only after an init

  P_SAMP : process (CLK, RST) is
  begin

    if (RST = '1') then
      rom_start_addr_samp <= 0;
      rom_offset_samp     <= 0;
    elsif (CLK'event and CLK = '1') then
      if (INIT = '1') then
        rom_start_addr_samp <= VTRACE_ROM_START_INDX;
        if (VTRACE_ROM_SAMPLES > 0) then
          rom_offset_samp <= VTRACE_ROM_SAMPLES - 1;
        else
          rom_offset_samp <= 0;
        end if;
      end if;
    end if;

  end process P_SAMP;

  --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
  -- Calculate rom address, and on overflow start from beginning

  P_ROM_RADDR : process (CLK, RST) is
  begin

    if (RST = '1') then
      rom_raddr_s  <= 0;
      rst_emu_gate <= '0';
    elsif (CLK'event and CLK = '1') then
      rst_emu_gate <= '1';

      --remove tc counter
      if (EN = '1' AND prescaler_cnt_tc = '1') then
        if (rom_raddr_s = rom_start_addr_samp + rom_offset_samp) then
          rom_raddr_s <= rom_start_addr_samp;
        else
          if (rom_raddr_s = VTRACE_ROM_NUM_ELEMENTS - 1) then
            rom_raddr_s <= 0;
          else
            rom_raddr_s <= rom_raddr_s + 1;
          end if;
        end if;
      end if;

      if (INIT = '1') then
        rom_raddr_s <= VTRACE_ROM_START_INDX;
        --rst_emu_gate <= rst_emu_s;
      end if;
    end if;

  end process P_ROM_RADDR;

end architecture BEHAVIORAL;

--------------------------------------------------------------------------------
