--------------------------------------------------------------------------------
-- Engineer:  Luca Caronti    [luca.caronti@studenti.unit.it]
--            Simone Ruffini  [simone.ruffini@tutanota.com]
--
-- Create Date:   05/17/2020 03:21:54 PM
-- Design Name:  
-- Module Name:   INT_EMU - Behavioral
-- Project Name:  NORM
-- Description:   Intermittency emulation core.
--                This entity generates a signal (RST_EMU) used by the test platform
--                as a reset signal. This is generated by comparing a voltage sample
--                to a voltage level selected as the reset threshold. 
--
-- Revision:
-- Revision 00 - Luca Caronti
-- * file created
-- Revision 01 - Simone Ruffini
-- * refactoring and generalizatin of the component (input rom is outside of the entity)
-- Additional Comments:
--
--------------------------------------------------------------------------------

----------------------------- PACKAGES/LIBRARIES -------------------------------
library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.NUMERIC_STD.all;

  -- User libraries
  use work.NORM_PKG.all;

----------------------------- ENTITY -------------------------------------------
entity INT_EMU is
  generic (
    ROMADDR_W           : natural; -- ROM address bit width
    ROMDOUT_W           : natural  -- ROM dout bit widht
  );
  port (
    CLK                 : in    std_logic;                                                     -- Clock signal
    RST                 : in    std_logic;                                                     -- Positive reset
    EN                  : in    std_logic;                                                     -- Enable core
    INIT                : in    std_logic;                                                     -- Init core
    RST_EMU             : out   std_logic;                                                     -- Emulated positive reset
    THRESH_STAT         : out   std_logic_vector(C_INT_EMU_NUM_THRESH - 1 downto 0);           -- Thresholds statuses
    THRESH_VALUES       : in    intermittency_arr_int_type(C_INT_EMU_NUM_THRESH - 1 downto 0); -- Thresholds values
    RST_EMU_THRESH_INDX : in    natural range 0 to C_INT_EMU_NUM_THRESH - 1;                   -- Index of threshold used for RST_EMU
    ROM_START_ADDR      : in    std_logic_vector(ROMADDR_W - 1 downto 0);                      -- ROM start address for sampling
    ROM_OFFSET          : in    natural range 0 to (2 ** ROMADDR_W - 1);                       -- ROM last sample, offset from ROM_START_ADDR
    ROM_ADDR            : out   std_logic_vector(ROMADDR_W - 1 downto 0);                      -- ROM address
    ROM_DOUT            : in    std_logic_vector(ROMDOUT_W - 1 downto 0)                       -- ROM dout
  );
end entity INT_EMU;

----------------------------- ARCHITECTURE -------------------------------------
architecture BEHAVIORAL of INT_EMU is

  --########################### CONSTANTS 1 ####################################

  --########################### TYPES ##########################################

  --########################### FUNCTIONS ######################################

  --########################### CONSTANTS 2 ####################################

  --########################### SIGNALS ########################################
  signal rom_start_addr_samp  : std_logic_vector(ROMADDR_W - 1 downto 0);
  signal rom_offset_samp      : natural range 0 to (2 ** ROMADDR_W - 1);
  signal prescaler_clk        : std_logic; -- clock after prescaling
  signal cnt_value            : natural range 0 to (2 ** ROMADDR_W - 1);
  signal init_s               : std_logic;
  signal output_comparator    : std_logic_vector(C_INT_EMU_NUM_THRESH - 1 downto 0);

  --########################### ARCHITECTURE BEGIN #############################

begin

  --########################### ENTITY DEFINITION ##############################

  U_PRESCALER : entity work.prescaler
    generic map (
      VALUE => C_INT_EMU_SAMPLES_PRESCALER
    )
    port map (
      CLK           => CLK,
      PRESCALER_CLK => prescaler_clk
    );

  U_TRACE_CNT : entity work.var_cnt
    generic map (
      MAX         => (2** ROMADDR_W - 1),
      INIT_VALUE  => 0,
      INCREASE_BY => 1
    )
    port map (
      CLK       => prescaler_clk,
      RST       => RST,
      INIT      => init_s,
      CE        => EN,
      TC        => open,
      END_VALUE => ROM_OFFSET,
      VALUE     => cnt_value
    );

  --########################## OUTPUT PORTS WIRING #############################

  COMPARATOR_GENERATOR : for i in C_INT_EMU_NUM_THRESH - 1  downto 0 generate
    output_comparator(i) <= '0' when unsigned(ROM_DOUT) > THRESH_VALUES(i) else
                            '1';
  end generate COMPARATOR_GENERATOR;

  RESET_EMULATOR <= output_comparator(RST_EMU_THRESH_INDX);

  THRESH_STAT <= output_comparator;

  ROM_ADDR <= to_integer(unsigned(cnt_value) + unsigned(rom_start_addr_samp));

  --########################## PROCESSES #######################################

  P_SAMP : process (CLK, RST) is
  begin

    if (RST = '1') then
      rom_start_addr_samp <= (others => '0');
      init_s              <= '0';
    elsif (CLK'event and CLK = '1') then
      if (INIT = '1') then
        init_s              <= '1';
        rom_start_addr_samp <= ROM_START_ADDR;
      end if;
    end if;

  end process P_SAMP;

end architecture BEHAVIORAL;
--------------------------------------------------------------------------------