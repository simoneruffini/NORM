----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/17/2020 03:56:37 PM
-- Design Name: 
-- Module Name: trace_ROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity trace_ROM is
    generic(
        NUM_ELEMNTS_ROM : integer;
        MAX_VAL         : integer
    );
    port(	
	   	clk       : in	std_logic;
		addr      : in	integer range 0 to NUM_ELEMNTS_ROM - 1;
		data_out  : out	integer range 0 to MAX_VAL
    );
end trace_ROM;

architecture Behavioral of trace_ROM is
    type rom_type is array (0 to NUM_ELEMNTS_ROM - 1) of integer range 0 to  MAX_VAL;
    signal ROM: rom_type := (
    -- put here you voltage trace values, separated by a comma (the last one without)
    -- the NUMBER OF ELEMENTS inside this rom MUST BE NUM_ELEMENTS_ROM
        0,
        170,
        186,
        225,
        317,
        320,
        348,
        413,
        403,
        379,
        369,
        359,
        350,
        342,
        335,
        329,
        326,
        321,
        313,
        321,
        329,
        338,
        406,
        472,
        461,
        448,
        429,
        407,
        394,
        381,
        370,
        359,
        400,
        429,
        415,
        400,
        371,
        351,
        334,
        322,
        312,
        305,
        298,
        293,
        278,
        289,
        299,
        307,
        311,
        314,
        313,
        309,
        303,
        284,
        268,
        253,
        240,
        230,
        221,
        213,
        207,
        215,
        222,
        228,
        222,
        219,
        218,
        218,
        217,
        215,
        213,
        201,
        193,
        186,
        179,
        175,
        172,
        172,
        175,
        208,
        215,
        210,
        202,
        198,
        199,
        201,
        203,
        232,
        265,
        256,
        245,
        234,
        223,
        211,
        210,
        236,
        230,
        221,
        239,
        253,
        265,
        273,
        280,
        287,
        294,
        300,
        281,
        269,
        262,
        258,
        255,
        251,
        246,
        242,
        237,
        238,
        248,
        256,
        261,
        262,
        263,
        266,
        268,
        258,
        283,
        305,
        323,
        335,
        341,
        343,
        340,
        336,
        314,
        293,
        274,
        257,
        241,
        227,
        216,
        206,
        216,
        241,
        265,
        266,
        269,
        271,
        275,
        279,
        284,
        289,
        276,
        273,
        272,
        271,
        270,
        270,
        272,
        272,
        266,
        253,
        246,
        240,
        264,
        285,
        296,
        307,
        293,
        277,
        287,
        312,
        333,
        351,
        364,
        371,
        371,
        364,
        343,
        318,
        293,
        271,
        257,
        253,
        260,
        278,
        308,
        309,
        346,
        381,
        422,
        464,
        504,
        541,
        574,
        602,
        589,
        616,
        642,
        670,
        700,
        731,
        763,
        791,
        817,
        799,
        820,
        829,
        837,
        846,
        853,
        861,
        871,
        863,
        871,
        912,
        938,
        965,
        988,
        1011,
        1034,
        1055,
        1042,
        1063,
        1104,
        1134,
        1162,
        1191,
        1218,
        1241,
        1260,
        1274,
        1273,
        1266,
        1262,
        1258,
        1257,
        1255,
        1258,
        1262,
        1273,
        1276,
        1279,
        1282,
        1285,
        1287,
        1290,
        1292,
        1337,
        1355,
        1371,
        1384,
        1403,
        1416,
        1424,
        1431,
        1419,
        1390,
        1353,
        1321,
        1291,
        1267,
        1246,
        1229,
        1217,
        1330,
        1521,
        1473,
        1436,
        1405,
        1376,
        1353,
        1560,
        1606,
        1638,
        1633,
        1643,
        1977,
        2041,
        1988,
        1947,
        1912,
        1886,
        1861,
        1826,
        1796,
        1769,
        1745,
        1729,
        1716,
        1705,
        1719,
        1704,
        1688,
        1676,
        1667,
        1741,
        2098,
        2066,
        1949,
        1930,
        1879,
        1837,
        1800,
        1766,
        1817,
        2147,
        2106,
        1972,
        1973,
        1941,
        1911,
        1884,
        1860,
        1838,
        1820,
        1804,
        1713,
        1725,
        1705,
        1689,
        1675,
        1661,
        1650,
        1639,
        1629,
        1543,
        1518,
        1479,
        1446,
        1415,
        1388,
        1364,
        1340,
        1320,
        1299,
        1350,
        1378,
        1403,
        1424,
        1444,
        1462,
        1481,
        1477,
        1466,
        1517,
        1550,
        1575,
        1599,
        1623,
        1649,
        1669,
        1643,
        1613,
        1614,
        1615,
        1618,
        1622,
        1628,
        1946,
        2078,
        1987,
        1955,
        1948,
        1937,
        1927,
        1921,
        1918,
        1910,
        1900,
        1829,
        1797,
        1765,
        1737,
        1711,
        1687,
        1664,
        1641,
        1621,
        1541,
        1593,
        1614,
        1630,
        1644,
        1652,
        1660,
        1668,
        1675,
        1602,
        1669,
        1690,
        1707,
        1721,
        1733,
        1742,
        1748,
        1753,
        1680,
        1698,
        1685,
        1677,
        1669,
        1663,
        1657,
        1648,
        1639,
        1580,
        1619,
        1625,
        1633,
        1640,
        1645,
        1650,
        1654,
        1658,
        1605,
        1642,
        1652,
        1659,
        1665,
        1671,
        1677,
        1686,
        1683,
        1625,
        1633,
        1634,
        1634,
        1631,
        1635,
        1639,
        1949,
        2134,
        2012,
        1964,
        1920,
        1878,
        1842,
        1818,
        1793,
        1768,
        1712,
        1705,
        1747,
        1791,
        1832,
        1868,
        1900,
        1930,
        1960,
        1891,
        1980,
        2048,
        2103,
        2152,
        2198,
        2237,
        2274,
        2306,
        2218,
        2629,
        2715,
        3024,
        3120,
        3303,
        3497,
        3482,
        3725,
        3438,
        3340,
        3208,
        3090,
        2984,
        2890,
        2807,
        2733,
        2666,
        2516,
        2448,
        2384,
        2328,
        2279,
        2234,
        2197,
        2163,
        2129,
        2067,
        2106,
        2113,
        2117,
        2120,
        2121,
        2125,
        2131,
        2115,
        2060,
        2469,
        2512,
        2829,
        2989,
        3066,
        3260,
        3239,
        3451,
        3297,
        3145,
        3022,
        2914,
        2815,
        2726,
        2646,
        2577,
        2433,
        2391,
        2354,
        2318,
        2286,
        2259,
        2237,
        2217,
        2199,
        2098,
        2086,
        2073,
        2061,
        2049,
        2036,
        2026,
        2016,
        2006,
        1948,
        1982,
        2079,
        2580,
        2560,
        2493,
        2435,
        2384,
        2339,
        2237,
        2245,
        2221,
        2198,
        2183,
        2172,
        2157,
        2153,
        2133,
        2072,
        2100,
        2104,
        2108,
        2111,
        2118,
        2129,
        2138,
        2095,
        2173,
        2668,
        2702,
        3075,
        3243,
        3329,
        3580,
        3518,
        3670,
        3807,
        3662,
        3472,
        3316,
        3180,
        3065,
        2972,
        2892,
        2779,
        2674,
        2615,
        2555,
        2502,
        2459,
        2424,
        2391,
        2361,
        2277,
        2239,
        2209,
        2177,
        2154,
        2135,
        2117,
        2097,
        2078,
        1991,
        2001,
        2038,
        2063,
        2080,
        2097,
        2109,
        2121,
        2130,
        2038,
        2060,
        2076,
        2089,
        2100,
        2216,
        2781,
        2772,
        2698,
        2542,
        2490,
        2437,
        2394,
        2358,
        2325,
        2297,
        2268,
        2246,
        2207,
        2819,
        3063,
        3358,
        3746,
        3736,
        4175,
        4090,
        4270,
        4284,
        4262,
        4399,
        4398,
        4466,
        4508,
        4510,
        4593,
        4302,
        4329,
        4237,
        3934,
        3688,
        3483,
        3306,
        3155,
        3024,
        2842,
        2790,
        2738,
        2691,
        2646,
        2610,
        2579,
        2549,
        2525,
        2488,
        2447,
        2415,
        2378,
        2346,
        2317,
        2291,
        2264,
        2248,
        2234,
        2221,
        2217,
        2212,
        2206,
        2198,
        2185,
        2166,
        2136,
        2111,
        2091,
        2071,
        2052,
        2037,
        2026,
        2021,
        2433,
        2718,
        2995,
        3198,
        3416,
        3724,
        3707,
        4104,
        4053,
        3786,
        3968,
        3978,
        4081,
        4317,
        4050,
        3783,
        3551,
        3355,
        3188,
        3050,
        2930,
        3184,
        3274,
        3107,
        2975,
        2891,
        2814,
        2746,
        2685,
        2629,
        2580,
        2537,
        2503,
        2875,
        3490,
        3515,
        4032,
        4100,
        4362,
        4664,
        4549,
        4568,
        4750,
        4615,
        4997,
        4790,
        5074,
        5094,
        5039,
        5252,
        4976,
        4606,
        4287,
        4024,
        3812,
        3631,
        3474,
        3334,
        3143,
        3009,
        2917,
        2838,
        2764,
        2696,
        2634,
        2579,
        2529,
        2398,
        2765,
        2950,
        3224,
        3552,
        3529,
        3856,
        3758,
        4050,
        3763,
        3962,
        4332,
        4240,
        4652,
        4524,
        4756,
        4738,
        4783,
        4701,
        4581,
        4235,
        3958,
        3724,
        3526,
        3354,
        3207,
        3076,
        2883,
        3209,
        3328,
        3535,
        3662,
        3741,
        3819,
        3876,
        3914,
        3597,
        3430,
        3292,
        3177,
        3081,
        3008,
        2950,
        2898,
        2784,
        2819,
        3224,
        3225,
        3441,
        3567,
        3581,
        3820,
        3699,
        3779,
        3915,
        3722,
        3554,
        3419,
        3301,
        3198,
        3106,
        3027,
        2865,
        2844,
        2858,
        2862,
        2864,
        2867,
        2869,
        2869,
        2870,
        2720,
        3094,
        3359,
        3447,
        3827,
        3725,
        4034,
        4177,
        4075,
        4038,
        4402,
        4513,
        4166,
        4193,
        4240,
        3935,
        3686,
        3435,
        3249,
        3145,
        3059,
        2983,
        2915,
        2844,
        2781,
        2725,
        2579,
        2488,
        2408,
        2337,
        2269,
        2209,
        2155,
        2104,
        2060,
        1957,
        1922,
        1885,
        1853,
        1823,
        1796,
        1770,
        1748,
        1728,
        1689,
        1737,
        1776,
        1809,
        1839,
        1870,
        1900,
        1921,
        1880,
        1892,
        1917,
        1939,
        1955,
        1969,
        1974,
        1979,
        1983,
        1895,
        1831,
        1782,
        1736,
        1696,
        1661,
        1631,
        1604,
        1580,
        1532,
        1595,
        1647,
        1693,
        1731,
        1765,
        1796,
        1824,
        1844,
        1740,
        1700,
        1665,
        1634,
        1609,
        1589,
        1571,
        1553,
        1499,
        1508,
        1537,
        1564,
        1587,
        1604,
        1622,
        1634,
        1643,
        1573,
        1539,
        1510,
        1485,
        1464,
        1445,
        1429,
        1414,
        1401,
        1365,
        1428,
        1468,
        1504,
        1537,
        1564,
        1590,
        1613,
        1632,
        1577,
        1607,
        1632,
        1654,
        1675,
        1699,
        1717,
        1730,
        1689,
        1641,
        1636,
        1634,
        1633,
        1628,
        1626,
        1623,
        1621,
        1550,
        1587,
        1621,
        1650,
        1672,
        1693,
        1716,
        1737,
        1758,
        1715,
        1808,
        1877,
        1944,
        2008,
        2068,
        2125,
        2184,
        2235,
        2167,
        2220,
        2269,
        2316,
        2361,
        2410,
        2455,
        2490,
        2435,
        2349,
        2315,
        2291,
        2270,
        2247,
        2228,
        2210,
        2194,
        2095,
        2172,
        2235,
        2289,
        2335,
        2375,
        2413,
        2445,
        2474,
        2399,
        2492,
        2567,
        2632,
        2692,
        2739,
        2785,
        2830,
        2835,
        2716,
        2719,
        2722,
        2728,
        2735,
        2742,
        2744,
        2743,
        2640,
        2619,
        2655,
        2683,
        2701,
        2712,
        2723,
        2733,
        2739,
        2613,
        2641,
        2659,
        2678,
        2692,
        2702,
        2711,
        2716,
        2723,
        2606,
        2635,
        2661,
        2681,
        2700,
        2717,
        2739,
        2761,
        2726,
        2725,
        3127,
        3169,
        3478,
        3493,
        3750,
        3532,
        3349,
        3279,
        3508,
        3454,
        3271,
        3119,
        2990,
        2877,
        2776,
        2689,
        2574,
        2590,
        2605,
        2620,
        2632,
        2644,
        2658,
        2673,
        2636,
        2536,
        2532,
        2528,
        2531,
        2533,
        2529,
        2522,
        2518,
        2493,
        2444,
        2404,
        2369,
        2338,
        2313,
        2297,
        2279,
        2260,
        2250,
        2241,
        2233,
        2225,
        2218,
        2213,
        2208,
        2211,
        2267,
        2319,
        2362,
        2396,
        2428,
        2452,
        2473,
        2491,
        2456,
        2395,
        2342,
        2303,
        2271,
        2238,
        2206,
        2181,
        2199,
        2686,
        2751,
        2649,
        2564,
        2492,
        2429,
        2370,
        2318,
        2347,
        2390,
        2896,
        3383,
        3281,
        3203,
        3136,
        3085,
        3533,
        3762,
        3576,
        3426,
        3293,
        3182,
        3083,
        2998,
        3014,
        3471,
        3455,
        3875,
        3816,
        4120,
        4152,
        4262,
        4256,
        3997,
        4284,
        4160,
        4412,
        4275,
        4532,
        4366,
        4585,
        4265,
        4401,
        4548,
        4261,
        4025,
        3827,
        3658,
        3514,
        3391,
        3175,
        3080,
        2992,
        2915,
        2847,
        2787,
        2734,
        2685,
        2642,
        2503,
        2455,
        2408,
        2364,
        2327,
        2290,
        2263,
        2239,
        2195,
        2118,
        2119,
        2115,
        2116,
        2119,
        2120,
        2117,
        2114,
        2035,
        2099,
        2196,
        2281,
        2348,
        2405,
        2455,
        2499,
        2538,
        2424,
        2384,
        2346,
        2313,
        2286,
        2258,
        2236,
        2216,
        2199,
        2142,
        2247,
        2336,
        2412,
        2478,
        2536,
        2597,
        2650,
        2643,
        2658,
        3084,
        3145,
        3482,
        3510,
        3843,
        3793,
        4106,
        3791,
        3643,
        3515,
        3407,
        3398,
        4018,
        3945,
        3768,
        3621,
        3396,
        3370,
        3323,
        3282,
        3247,
        3217,
        3187,
        3163,
        3140,
        3013,
        3472,
        3463,
        3877,
        3809,
        4150,
        4044,
        4336,
        4059,
        3839,
        3684,
        3551,
        3436,
        3338,
        3250,
        3173,
        3106,
        2940,
        2948,
        2946,
        2944,
        2940,
        2935,
        2932,
        2932,
        2928,
        2763,
        2694,
        2622,
        2556,
        2499,
        2448,
        2404,
        2373,
        2314,
        2221,
        2193,
        2164,
        2140,
        2124,
        2106,
        2087,
        2067,
        1987,
        2033,
        2116,
        2187,
        2243,
        2293,
        2337,
        2375,
        2405,
        2312,
        2386,
        2446,
        2495,
        2539,
        2576,
        2607,
        2635,
        2658,
        2512,
        2528,
        2984,
        3014,
        3420,
        3385,
        3719,
        3648,
        3919,
        3772,
        3667,
        3580,
        3501,
        3427,
        3362,
        3310,
        3267,
        3075,
        2955,
        2848,
        2755,
        2671,
        2597,
        2534,
        2478,
        2425,
        2332,
        2375,
        2405,
        2431,
        2451,
        2471,
        2488,
        2510,
        2503,
        2365,
        2320,
        2280,
        2247,
        2223,
        2202,
        2180,
        2158,
        2072,
        2123,
        2211,
        2293,
        2356,
        2416,
        2461,
        2499,
        2535,
        2429,
        2432,
        2433,
        2431,
        2428,
        2426,
        2423,
        2418,
        2415,
        2291,
        2262,
        2229,
        2196,
        2168,
        2142,
        2120,
        2108,
        2071,
        2060,
        2138,
        2197,
        2248,
        2300,
        2795,
        3225,
        3148,
        3045,
        2924,
        2912,
        2902,
        2899,
        2904,
        2908,
        2907,
        2907,
        2791,
        2771,
        2791,
        2799,
        2802,
        2800,
        2797,
        2793,
        2791,
        2643,
        2572,
        2506,
        2444,
        2387,
        2335,
        2292,
        2254,
        2222,
        2140,
        2178,
        2203,
        2219,
        2222,
        2219,
        2216,
        2213,
        2163,
        2103,
        2119,
        2129,
        2137,
        2139,
        2132,
        2124,
        2115,
        2023,
        2028,
        2052,
        2065,
        2071,
        2075,
        2078,
        2079,
        2076,
        1974,
        1956,
        1938,
        1923,
        1910,
        1899,
        1893,
        1884,
        1878,
        1806,
        1815,
        1817,
        1821,
        1825,
        1833,
        1848,
        1866,
        1840,
        1835,
        1898,
        1955,
        2010,
        2057,
        2092,
        2126,
        2152,
        2072,
        2003,
        1955,
        1908,
        1869,
        1833,
        1803,
        1776,
        1751,
        1671,
        1665,
        1656,
        1650,
        1643,
        1635,
        1629,
        1624,
        1621,
        1590,
        1665,
        1727,
        1781,
        1829,
        1872,
        1916,
        1953,
        1943,
        1889,
        1905,
        1919,
        1938,
        1953,
        1964,
        1971,
        1977,
        1964,
        1934,
        1907,
        1884,
        1862,
        1845,
        1836,
        1827,
        1816,
        1811,
        1807,
        1803,
        1798,
        1796,
        1792,
        1788,
        1788,
        1837,
        1884,
        1915,
        1942,
        1968,
        1988,
        2007,
        2023,
        1988,
        1934,
        1886,
        1849,
        1816,
        1786,
        1756,
        1746,
        2066,
        2152,
        2078,
        2016,
        1963,
        1915,
        1876,
        1839,
        1806,
        1832,
        1870,
        1907,
        1933,
        1953,
        1969,
        1984,
        1995,
        1991,
        1975,
        1963,
        1952,
        1950,
        1947,
        1944,
        1938,
        1916,
        1870,
        1831,
        1794,
        1762,
        1734,
        1709,
        1688,
        1662,
        1594,
        1587,
        1581,
        1576,
        1570,
        1569,
        1567,
        1563,
        1519,
        1526,
        1571,
        1614,
        1651,
        1679,
        1703,
        1726,
        1747,
        1676,
        1687
    );
begin
    
    
    get_data:process (clk) is
	begin
		if rising_edge(clk) then
			data_out <= ROM(addr);	--get the address read it as unsigned and convert to integer to get the value from ROM(integer)
		end if;
	end process;

end Behavioral;
