----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/14/2020 05:43:53 PM
-- Design Name: 
-- Module Name: NVME_FRAMEWORK_PACKAGE - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

use IEEE.MATH_REAL.ALL; --for log2 and ceil

use work.COMMON_PACKAGE.all;

package NVME_FRAMEWORK_PACKAGE is
    constant NUM_PWR_STATES                     : integer := 3;
    constant PWR_CONSUMPTION_ROM_BITS           : integer := 10;
    constant PWR_APPROX_COUNTER_NUM_BITS        : integer := 31;
    constant INTERMITTENCY_NUM_ELEMNTS_ROM      : integer := 1000;
    constant INTERMITTENCY_MAX_VAL_ROM_TRACE    : integer := 330;
    constant INTERMITTENCY_PRESCALER            : integer := 16;
    constant INTERMITTENCY_NUM_THRESHOLDS       : integer := 2;

    constant NV_REG_WIDTH                       : INTEGER := 16;
    constant FRAM_MAX_DELAY_NS                  : INTEGER := MASTER_CLK_PERIOD_NS *4;
    constant nv_reg_addr_width_bit              : INTEGER := integer(ceil(log2(real(NV_REG_WIDTH))));

end package NVME_FRAMEWORK_PACKAGE;
