`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kylT7SNcZwYZgnvMV/JDafym6dB1mBLeeUv9XKg0HfyqT8CXaBGpQFOQEn5SUK5kjlX7ig9yv3aB
8QwHm79ZEA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nRmypjT5263UN0z2JRGN68ZwlwA03XA02rv4qCb50yJDmeb6PUU/EJiNMJKwif4h3vH5woeOWeRy
AijHIuqOfQ4Y7t2rBAoEPGKuOXAn+UMx9GWMjvN6BbLKUUAvJbiOVRIwNzfSPiXJ1lgqf2O3eW/b
ogeX12/EsZTmuHhflfg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bn3LSHWaAaOc9CPg3uqB03bUA1MWUiMLXiUYc1tcYeORvB3ZCgSFmuoBCe26FlDNSwtnn0Jqxifz
o3btBDOb0Mmvosha92DoVWHwxB6gi/QrpkvxknAO48sZft6jmY8CAJytKfh7RzrHUWZuWWJ1KgWo
hy1dGyGjW2+08sKMyc6hz1W/yOA5r2GfXsXh33yV9lpFSQVi8Wk4vt5+LZGLws9zbdO0KkTptOn6
0u852C6fGsbFA/pFUAwcMGtdDDMuV0I99VTSlzQ9hCWfuOmrrQ0nsujWSG9jjO0qFFU41BP3eHaI
+laJUDyi30VecEicRBc/TZrZ2QgbmDC4+wqgow==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TqOIcExxHAhmDTmpMT3XPkBmPmxIqDA0+ljPx20AefdYG5wvQKZ69EUD71vUIuMoiTW7aBWFb6iw
TerEWkf2lQV3TFPkD5JGhJYQfxj+KC2j5S6Ach2MowAnVSD9M1UPGVAurW5lyUPG3fpAVOSFTMEI
1fJ2jNmKjbyV0X7zdBTty3EceLk5rPe/ADw8I61vh6Pd7Rf2DiZxp1cpDzRYvsjoto65wAHpehwG
yPVog+HIsZ6UlcdWZA87FLyK6QCycalPe19t2u869YLUw8tdLjCilZqTNQtDqSEkjqZe7D02RW7r
HnREQ9tX3Mib7Id2reHfTnxITPgEjiXNydI6Dg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SmETBvyvplz2+YipL8ciNdINvEtlNK7HFUk/REbiiPAvXSg2olq/+eJtvzZXSmQivoPOYj3MNrtd
DORvY6eVr6kS7hDmEl25ZFhVAepL5TnAHy44G3d/Ffl8Lj+hMICAmNZTjHhxm0SK4dHfwv2GDGHj
AgzWwhoSMvp4fWbDR+MouAkH+GL9VflGzzwSwk4iacctH6GMBWkJFjxG4bD1RbWVVMjxx4FJ2NAF
Wn8BCAi8a83yknuiBDnHUQXXKtA6BXnL7HRZy2Gsp9CZxRx2lKYkm82QMD8R+FqLsztFuDXNWSKl
awswsqDXhFO9A/2Ge7af5vmt1fhTbpaIPrusLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
StW9wDeopWYi8ygk17xZzVyhJcND5ccVGEPD3xxFtJPyhWRB9X3RnS9jSSxmyhC0ujqBzfu4ikJ4
/Eme6FW2b6TPVE7geg8soNIzuM1zCFotuvMhX5I55SDjHB5NR1kohZOEQmMXCvBjKMRVHXeBnPsh
c8BUoNnxxEYWLWpb0R8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dgt7h/HGpPE0xZc+ocdHKDopQjEYTuKgWjeOzNBMVcETRKCabsWXtyuBcYIsZvdx3mYGjmnajHsY
zOdzJ3SSVV7hnxRdS2zmQgRu63nC7p3Vn4jmWqF+x3OrZwEkmmV5NXfRAc0D2Wmj5ROON3Pi76L3
K2d3FDk88IFYU5GX4IbPnF/v4N42Ql6J+e7DMh8/ZMVCAMUl9FWeA5R3RItTY6dSQMF3zFMpxY9q
q7CINCjzdmeCGbT5fdIaBJKy8hZh19jITYg/jVRbZm/LRLpCxC2blt8IVaHB9G4Yr+rzlXUja7C+
BlJQnMQF+OTfORcOoLWElotSL8GEMVBes5F7+Q==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v6KS+vW0qRgTnr62oMcesnwexJfTvKFWjrSifMejJmZuvtmyHbptWIjtUMoFG0SqggklSdAV9uGM
XBeRBSvpnHy68h+I7eedV3cWubOxIPL8Ull1muXSb7YtfIGZipN3Nfuu9exnMxlHNC2tpzY0E6X8
UE/KoOhoS6ZfvS3P0dyyCwYlBTUwc8UbGQpVPXrPdOYuriyWxCibFzjhJzf8UqYi8OlDUV+hkaWw
535w0538ACN0vuxPz4WuvqYeslD3RM3X2D/XfMmEi4QXGNtr1BdZHU0d6dWKKCfzG3Q87cTUTgef
HIRoyx1ke+QB8TUpqmmmHX/wGTkSLhPPWHg72w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98368)
`protect data_block
n8DZCN9Vvq6qoayNtYRIt5fQ5smXfgNQrHXDdjByi7NtD3BjADAkHxXpNrCMdgJyPETBT02CY5an
6inzbRqx6BTMeIiVY7f7OxXtb63xFVgtn7/TmA63UrPKvx9GaAEGX+WBYliQf+/WkcBkU/UseJ5C
xl7MXEMNYOO1KneEiz2hPtTh01kvs/Q4OVVwafTm/QoVMp75ddz6z9uKG0FugWqd89QVF3OTh2Ue
LpbTx13pPhDkpFqYMMYNd8J7BDsmlXctT1jlvB4GiapLru1omh5a19kKHazt4dtUBIk7F/u+nh1p
1RSWJHL2pKFnYKYQVgfGO6uLAWREGu0i08H90VnkpNX3qpRKKNR4khI7b5N/lfGApRu5LElCVjnr
X5xOtcJVY93a0Sdx6wE9i63YGy3mkPsyLYltRBWWCH79hljp9s9AVz4mfzQ2aZzcwS+zY3FfzW1I
6VgocOybDywdIaHX2ue3lzEClcDgbxh103P+QBiL00VzVzlmgUeqQ44QRuvm1jgCmw/xfOOayLZL
ZzB1su58bENNkDgDK+bXdcwQlSEU3E+ayhsPwdfuSGT9BmvUNah8j0eXD9W2jKwOshkWmszYPK3g
BuVXJfJd09ykreAEGIta1c+dK7dNv3g8BaEVuj7eQya3PzDpHcm+WcyYhRItWRynjrYzxldUUm32
Q/Cwvjl/VFyOUFmn2qwB4wgr/jl3sCx+1bRFweie1hyRHeOk89hQQR6II+39zZB9qMVinWUTTVrA
ZCwht3sTZAaKYQqMuBD3EhjYktP/892xoLj/GegHksm4Vl/D0PaQMfvAR5U+WrXWSi2zxhUDJoAV
hypIQXzGl2IWaF+iFIV78a19GkwOkj6T6709HLXYB+/SVLG5e1RUgbKk5vRMTOIi97yCx6O08ImB
tkF7bFcat7gfUUG+SX8VcWazsFLGdTaRynMSCfgBbQ2Gu7tq6btxq5m9Q4nTJQieC0fm70WHZHWh
i+1k/1FWsTUA1HPVAQcNfVP3vY0IG4wY/z3E7g/vchBoe0HMzO0p67MTAsp52ESx+18WR43zDzRy
ZC9mwRY3FridUqj/ygxoFt8CK73t8RRYpKhDQFcAVZSrXgSpx4pJh7vQybB+fG6Sn5WVu39XGINj
FA/PAvy3WYMMyV3KUC8ZK8izl28ati6dxEdsPXR9z09c7nCR0vmSt2kRTkmzBdGzt49PoMIQhZnQ
HK4PgEmSXHrL3duMjtBSMILNkTadDEO4ofET4+5kr6OmUwpDGNbPGB7wP7I8aVxd4ZCBKtRcI+8r
8/1h7WYvE04CtGlLCIJCiZtK+3Wj4UTr+frrTsBf7tXnWTH0tLOeEWLTg5AClTapirh/f3qJlLPz
ik/Yiroh/CL4Ep/grfGncB5c6aSHfRUjL0KG5P7PjyA5NHVN9fby0YAfiz7yzrZNF6oq34k/HxIb
go6Yqti+TuxIjA9GqYnxzhLr+bNH7v57OZow5AmiQKqzOiBLHMUq689oGQsQllNg4WcEQoiQJBmX
AuHwpWMB8T6SNBuy/vL14538Vles2pYDjbr4G76KHy9vJQyKCshKGjwdrsAjapiv+/RFzFTewryQ
IINVPuKQxGIzbfrmKSRpMoMJGa9ZQGNpNes2eB+APDfFXfJpYJYTRUh59QR1Y9Lh5FiQfa8cgWhy
dJ7khaT7UK7nTrPCLSKVfkXPc9pMft1x+kuCSrr0+zWbl1FJEO5RNOMWBYiBDhCUwlxWRxounWgu
G+pIdXp8KIVUmS154jtPyaHVxa5Cg4fcS0TWuWw5D6TkLuiBXYRPhVWYc13q+zqdypKHl4F309Rf
YezWfmfUQb2HiwQVQ2JTzIp0Su3DHEf5RMd1RL/vYoDbwiECwHPGMe8zKrAQPT+x84dXoa6uSoGJ
cIyyhXxsyO4v+DQM4iH+5m6DqSuI3z0VCMQxXg9PmFwx5UB25AM7uWMtLjf8HZ3nECXXaGUPdStO
uLCrk9alyKasE02jLI75i7tdM45rOY9zbLmsOoeloJAfmK16mvKZi4Nxt10BXl29rxkfusGohw9x
YUIbbAtLiPr6SyYZmvLTum/5Jy/8Xa34kodBL0fOszROJ0I9WMiYF06nQrzVjl3E4vQFcT0T/KxY
ccCeEPKgAaDrdSTTLJFRVnqhttXU3Uphn8LF4voYhq+I8zp/HN3EncQX1U+HCa3qgoGl7GAKCiml
OOrYDxdC7zBEwvPS8ph8s+FmvKOzaDI00HG0HZ5HJcoDgFl5mB2VaIxk78Wm3+eQGymB1Pl7464O
5sv8oNzrwx3Oqwfr1FlJ6Jw7fyBeHI/R/AvoTnr+/2eVxR5SWKJ0owpDxl4ogZHunpcRAVN+JAKt
V3xe8SiH0sgp5EUAeW4a2amRoKIupfzJWXtzErZ9mW02szTvBfE+tT/6zw2c+mKfX7I90OfRkxMX
3fz4nDDO7EGdQAkDng5dRiO9BISf1266ll9S5WIvnfyzptmQZkz1nprAC6oSZyrKS65+J9FW4QnT
BUCIT5m9H9fbI8Zd+SWANMKbZaLUrJtsLPQ6pGoKurvllrc52g7tn12UQvNRDlIbuuBauS12b2q6
TsPLD/ALZ7ZNQdCFt3S7bVeLm6o5stCT5l35dsJbkssgA9n7JrtsjuX2ILOr44BrQT+fE3cXCxwJ
actbhUuN3Bhw+CqNS8lErMw0imDI6uFlbz+m4u/rA5nn4/LjkS/lALcfzzbZ/mUUwPPxm2hnqCo4
zK60jKiQNSjV1Vel5KYaP7N5Xz+g/jZBYrfHEAIQp7S00q5vl5gQwEdezOs0w1dIhVSs7ZczRGJQ
dcJhUodjnal60imNf1W0E6AYEr9bdRKSWO9x8xJmfinHeNwWYEm81J4dZXFHZR6lGyJ9lNE3RS9N
o5QFu7uN7KYFrnmY3mr+xrJoGFEdaEgDVpROUG1zqV44D7XyNHOedzIECV+eGMsdQqwpRPGY0sRs
9G2WaoMr7cogr/OYEslYFJY3RUUyZhSDfj8ck2/GAaALx3wvG+o1dTWOBoG//w1c/IQmWXUh+Vh/
Pax9i4v/CrNLwZx36swuEDIUjIzJaZ1pIeBQhIsTFSC5lvHW8D6jlQeP7fjSYKqFQY2KL3yrcNu+
Bj2ngCKN6oqvwEs3s+ophXLvzZOl8N9VL2iA8kfkgvT3EBtgVDdpEZ7vXRr2Uk1aUGH/gk6OCU20
WfLTEl3WNe30FbxOCcJFXyQTHCYotrmJw/Zz3jsxN7zCJiHulReYKTfFhZzFX23Apx60WYifZqoE
cmGY5Y5kxzu0ZXAEIZe9FoqH15l+vJzPFh6m7hXF2YlvXz+zizMpsJvZVH72gVvB+85z7xVWvnoh
L+tWoMD+YUHnCQE3nkTcj8eSapg7tnEwSD2zRgz9rASDjTEIdrt5bkIpU3J3iGvcsdqTT6uf0pf/
xh4QoBGQimYRR96MQIWpslmEaFs9H3tPJGBagpe8C0fraQOdpojrQP/3eEilLVkWI/I00fFePxo/
nb/SK5yIRrwCgzM06LCeY15CwbuwF4mCndwOHi11R9wGlERnXWpXlskwiUSZ4ll3MV8+V8SbWnZQ
bwloY6ss0vI4uHm9bVsaTCoM6Qu8f3Vmj28mDfd8ARJMI5thOGViGkpaqpaaMkAMRyFYbhSx3SBd
Y7mKqtrHj05aQnY3z2p6vsem2NKETUhatUa9yxwze65IVUYmHplUfrePtiQ0n9HZaPNoLr3rETZ2
yfCq+w7LYMvME21F1zgdJsSNkgN3613DXkjsTMcw74k5exZTqNd9yqTHwxQaiNPbijBK8zquX9pK
xD9ZxHzMzq8LbocfxKBtFfj93E4WZGhYsDGcxfUiqkdKXhKV6C6VeI+obwutWcOOU6BP9pmVuzby
7Rz2sGZzdPRFQYZjFGclVxVAudnV74ijF94b/6Lp/t3g08AwDcfA0Xtq/TQD0Ez7WpDQ8oDCzdzh
isgcqbSzXnXHn1Q9pA58cThQbBZk6e/RyMXxp1Qp4oXHnCUrOMB2OSFkE5F9gLXtUrnxPraT7fcC
fK35HklSEY2uIZmqXg82/mtG31u/QQvPJGDkM9FUPfmzqVKQXkbg1UBsbGGqK22xcUtFm1NeJmIb
p6N+My5Q0a45pm+dokGcIzHyBUgRXNileyLZdBZQK2qODfAqI5wL47Xb+T9GGOuWcN8aJaoUJn6H
RkMddhMinmKQ5WaFJPSIrA/Ul53bNdWCPNpnZKnqiAwkJuNe9UMfG1Gvn9R2YabEjRL/1zankKw4
dQrm9ebJhkvHvz5XV3xPk5++KX2X/r0YHgUeZLr051WTgBF9Bgtz5WfnDyDBBhRBrkklImHd1RQN
0du9yzzrTW8eFuYOsVwsHZQZqS+OvAZz5QTEB10dYNCrz6pR5WnL546368eACS7lfBOW9GNeeKYQ
+cLNwAcVtC05dLZTAe9e+d6OdKZw7uIJWSJNFfyBJJTutL4IlsBJSWBjyHokhPXGx6UjOrKvgcLQ
/wyHb5MksEJQB8MqWPVAJZkvapaowk9KWrnSNgvCIMxRcmQW3A+HROXVvpRy1Ra2LMJr2zvrZfg2
d0S03NVLsMjg4RRTlvI7qnBxE1oB4OCEjNB149194hrRCxFna8xRXlPr5xIMg42BjSO/LioSchUx
uGbAvWx/gTBBvnptmZ1s5Xi/fFu7wLWw8hzz71CGse4sRTpsyl5rntGYjVqey5LD9mpMWXi4KwRI
hNyXiIAJvr25Ark3F4MW4OJH/XfMB3M0y/QLMYzCBcmIcG4I0fY8hwEpae+Ly86LehmI5cwnw1Rx
mqbvZ17qtZsfLmhd/s134596P4xw6lgsnYftaselk5pXJy1jatkEEJhx3JWyXvVIqEWg+23jdriJ
qTxbx0whlncVwad3eFullDOPNPNLcffBmj5kj60rbaLVVnVUAve0neyrISl/dVHX+VYJ1U4FMUij
ykozU5NS8ulDqydakdKLVL1Nd8kjKJQ915fIPTkXCVfH4COYPErsdCsTPmGTs2aS+hBAatY6Yymn
dCfLSM6MeK84G8MNeWQ225viB8NbwaRvpW3tmHIXyKREPC/SwGjXXnyLIoh9H6kuKT5Wn4/ac53/
BjAuEfWo5qwnyfLal1KKpFvOIyYj3bXEfaKhbGbGGvdLsV2OxWPoanrqrbzIdfmNbEbWDExiBqL5
g4BjRAPLQ9YTS0WUp9bbS+oPeJSEcUZ62+h89PRMMpjIwm902fxHLfZg/BpVDoLDrxTtVZL5iT7a
xJpcSYKPeGFbG+SsMAss67np/1y6iOY4k71MRHK9D8VbRugBTKoCG/mY38Keqx5M43cswozIRhLE
K4LICz9SAjEOUQrwpAODC9Bc2V+fZcwGN4eCe6suJI5AqaoQL5ytoVJjt1qlAL0r1LAhXYFxPnN+
2ST5KzWaDpQ4PkEwW4kyXx15PlKIPrQGttwux8CUQ4S5mdqOaco0vGJWvnpioD9mi7pO1FkTKXvn
d9XUjfIJSUtfo9zpBctkS/AQTa5uYFNxUechCu5RZ0jWQNkx5Iz3cbP/WRqWMPMHy5uzdyb/NZGz
RtUeVIIteYuZJz69CRq9MowKAIGqJy2i8+MPtOlO4yMRQxNw78pQqqttxU8daThTAuw0mon+mrBn
THfzoRCAy/fadVf+ZpOvtPf/spnvja9An2QYhExSbKshmj/nAZdsVvc1Ek+jwEaVlkzsQ1gAcpDH
ZDIPr9PkoRqHDTfPciVfSw3i2ml8H1etSgfsBv4auiFpU28NPjvjSIHWGxlaPgAs4TfNNcNKhoJF
EsLDODzDLnz/FQaXnikgFkrboqsX/6MHufB3DbviNLh3x4bZEMY6wm/e2iebhojzTly6mlEScwec
laEUiCMqk/zp9Q7rmx0MCF343/7LFGHKwlgIckX664drPS/6C3br7NwRqSo6ga9f7o37sor3+A02
PHoUhq2UZy7B/11YtimMuWI/MeiohAujUnpPgYiA+AHsZd/mZHTTS03JtFtKpetq7wocGVtfoHJa
oKhr7i3ADmfpciSy6UnXjRKHDrSZttDvVgzJEoHXc2UexaBhRF1A54/FbkVzyN+fMjp4KWW0yAYF
/PMJLLDlc8ZNd6hWyULD1oA6X0nrRv4exR8MfWRwQ0xSmiRpqGRQmmNpvGHpg52jyG4Di1Nqh/8t
Gq+GnptivFO3syPmz//64NUXBAhCy1Ts8tcgFxwrF1Zi+bhVBX8KqsRc/tlEu7C3r5udh2qaAGo7
N8evnOPDs/CtNqT++JL2OGTdrWwQhCePaKtUgzRUnn7/ieWgsJcIBENIKiMTbvLIL3JJ+rjGsllB
NFNi/OZ2UJf8xSPulLpGdaXtNJR/DEHB1RP9TE7UnVtiwIYSA+ZEvzHRcoAWTKCxmYL2U0YpJ2+J
b0kAqfJlsnLObIIDIiJXW6X28V0LvFcoA62372XMfZ4OKOR4L7fZ5w65VgzKmcC8PH/TG1jHGxGh
jC2WFpKRxqNxvJNaSleCma1Fa6yGI04vpMP4IqB11nyMtDFt1asUzR4T3UyarM2dYpFRb4vsCvrw
lNvdmBBCZ30hW9ywTTOi8qOt5yREkzSRSi4TKFYnSyqkPUeCUqRD2y9J7mlaJHjPTMvmcWwgeMgd
v+uU99sTyy8Dn6WhDngQaUuoRA+SwYrwXL1vNOS3GSKuqzEa+CB2KSA8zQDa1IsMsQT/Pf3OvI6U
kxJ7EdhbEMR/8p8b1MvOPk10zuHSUmqJ8a8kQgs29Z9BidHC9ryDMUY2wUB9sz4IW7by1S12ffYx
v7+0e5i2B0J5wFV01FDw131XVUfWCepaGPWSpCgWLHE4Jsn6wS+QQhSIa05mXUza9buLpdEaKQpD
DAxGUPou/7Ygn0G/EteJl5Moqc4iO3+/qmV6Is01Xp3eoAUylB+FU/PYSBB02XNEKYxi7fAdBMIb
rdh9bESoS+xPTLKyUnI5uBNc8NK6o6Q4TRI492YobvUdsaqHhNkcER+BVsmdRKo7ELBqmZ7cXEN+
izsnStfZQJd9EsXCFYXibJHTfCfuqSwSNTGZl8UEw1pEsUCeEq/V3VQ53byz/bFT4A05gQ/A4tiO
Qw0NnbPexSlYf31hAoxtQvgi+GqyUUKyxCZociH3937HCHrPZ24zAr/0PEbEr++0Hm51A42FrBi0
ELlT0i6VhT1ei2i+s8CBAQSrqTD0x9iHZ6UQJRRXqo9dg4EO60xzKAh1/1YrP/LoZ0W+S/w3VRNo
OcssGSGnLNye3xLlPxgNy3LEh9FELZcdFPPQ5vPf/L7LeU7pv36ZWJ//6sjTniWK0LXJa8z6MFjd
Fvx2WtOx6vKwWJUnhIms+AcZmlkX9rqVTDAZq18K0YiEpPw9uGYit3ziM3VLXoxS1Rwvw16Pie8S
1I8AA3W5OdmBO5HBOlG2mbTAipcYvHswlBGAdrQ1hT1UMiRry+Ru8bohK6HKOY895W0YiH6s6qZg
60elxuAAdGqWwGE7K+CxCOaH3igkxryvLlQMDboSRElRjHDE+TUPTfr7TLudCsIUgJ59i9ZfRNd1
mAgryHxdyM1LIOpRcc7G4it2fpMJW21AsWZSFjNio9xO8rC/MAzjBIkhJVNilMSkh2StZpyaciJV
+vEXTGQhUfOmiBz/Cypbjd94osJgQGRtfS1tpV9Dz7I8O6BBt2Az7RR5UbeLs/lj+oZIRzL9A7tv
QHNgylXib0mRLVxyPj7qILgkRYTSN0EcJZ4E/Z8mtXF1jHCK4W1/KkhmyxhvV/Endd2Na4g6B6a8
SWa22ZiqpnfRw8c3fjVpTpvF5q2VqRzSqHh+uoeJvLg2HOnGzNWrFn8JjzuIm6i853pqG95js6EP
waI8yWp2AFSpY0Y5JPC+XM8MRoG3si6RG+PZPmpEpgKyWtzEPDv0jQA4ZZGLwOi9anX7I8IO3z+u
fSFePNd2nGrl+9FnrzlHYtqBZZtQU+8S+6lIW8x0peay/lPawYi+uDsAifAEmKR6GULOV9f+mVNH
677+6ZjamNuGokrBaEWjEFLWnnv6FvoZXD2s96WjQibeXRmEWDeCA+bMlGX+6qSRroFJHqzcFqfv
lqwfV8L5qcY1evp/ptO/g9s5ucrQCRpec0uWpW0Kuyia/Yl2iDLmr5tmhL1TkONljQJuKrlzGl9K
H9scR/1y/yVt0dp8Yud0GtpUWexuQbZY/RyECbUk7FwDo5/dgsdK2NDwpsYTL1YSr6JmQjdTLJkT
yP+TzSFM4Iuav62s2d100v3XRMKwM5WD8bfmuZBUGtJZTHTHGziaQuOv/uHxEufD/zJ+YfXZF5Xz
c51BWiAJwn5/rQDMRW/CIYyotzPMUoMx0mSaX4W1qAVoPfXffNfI4yFb2FfXLj7g9O4SQL5s869m
xUoPWi3iIpHRb1ADk8EMY7xAzOBjc0NI5/2GEQ+iaFHDEcpxUEnHDUmZQXFgy+Cf2ikjzVGr2x6v
DZ0FV14XsKCrYeiTS9A0Tqc4eON5lBIn9piTedMidcJHAkLOjZzon7L+mb1gZIAUBUoR/o8wBnMx
+3OouFZDCuWUofNY7WGQVhQfE6iBwvKo1bMEiqSeZi8s5CqtZifqcWJ+8dpJ1jwxtTFT29hcfRF5
3nfyK89oZ6uZqcr4mqJ18SaAwwXbwPFFEZ3tAXhU8k2t+krba+Ste/SEFhQ0jBdaW7uFYHAXXZ/1
l1f/K1Oh/rIKb/d9gUNMLsdIYUCdC/JJ1lNPGWRj1lmebvXHfzgYg3Yw9AsWA0u7+EJWFTrI85hV
mDjd6WqRaNGWE2eVGHtEbFkejmzmhv8FFroLcXVoO7je3NqpTbi82cBylqj+XjYmsMPs0/r6h9Gu
5JnPfkznV5wbMwH48nilJkCkPmtYXFMuPws4OCTdpLTPMiBoLZTYHp8/rXFAD3lQnTHtyzMNZTzG
BdDeK1UyPRx+dZrj44GxEVb179cI9SzSmRMPmSDHBKa4pTvpWzoXDhUML4TzwgF1RnQwhYpgACgb
ZdNGoM23EcK72NOsEN9LrgQATlgK/6L38lRJbSaEslcC+EIcsr9c4hOg/56ObhCCQqIcmS5qWQfG
vwmHnR19htDUvoGPQnZ8W9TJiGWPQ/MoB6FJdcsplC9kuBzZnv07g2AKct1Uojeo9I9Fu1zGm3pp
+MSHiz83hg4pd3YOnD6lr3YCH5/2Nh+lptOs48ZdCp7ApD5eqzROR+0yFko79BL2CHufelCwUOgV
gyA5L7RhvdmSNPa/rtWQ6P6sUQt+bzK2jUVs6skTtSIMLUGiwO+AT2O1S8pc+BOvrhoEBiZeBoJs
oP6JjlocX/i+ULZadYJT7XMwSx09aj4w96LPB5LRo+fdmOSqJfz5GYGFi7C64P8CFnEZ3TcfneeQ
rPUnThkKwIv1fTU2yLvBMDM0gowaKVbXfVp2hevCfUubNOQZbWJHaBgfmcPrEHXg2fH2uNsx3KWO
KpUYvyx4/GlBNXlul4rFv6Oig2WaJXXbiC9lfQ1Li497O3XoLHfE+yINg1ck31lpEzauUOFIGR8j
fk4HNB16nyLc2rZHvHwV9BT4KavZ2acJ/YqOqcPQEnfA0UC25vN0iETLGie5jiEdZcWdGwFzW2rD
WVc87877HfobFf/bBcSLjg8xZr7MYj9mlYbbFNu3WbSlPlV98oBzDQdvbSmn+vaTyI1ykL9bsew1
qYidZYIVQrY9PteDnzYLuOyEfomABKtdXKAAf8W22iOleMBuCr6oCWVsP/IbubKxx95A56tkG9c+
uv7hs/CPwpav0ZpvkI6N4U8xRUyuitHMatffrg1vyRnLdSQsXsX6TyEyr3TAmthzggL5OS984E88
OEW7nTvsfOIKh9vKm8KB4WsTUViKCLbGay4lFuOn0rYdu5mx1d3/ZX4vGjVimNTWNVrhXPFV0A/j
UfHFY7KpF+3ZQAeFqW03o0Z/KRVN5lyrJFqg+ZBBLBeA/98P5LjbyM/fG9ixEsW+1epgPXVvlsgI
lpKbCoJ5VEDJ9uLIyz0J5yIxXIxmMYMG5mEd0EVCaoH2gaVL5yCd4sCBYpLApYRrXXrtIN91HPix
n+jHh9GGBhu0mGofTmfR0qFsFAD77tjDf7hWnefGcTqaBSZVbrr3JbZKsxPaPbfApA7r0KtLSXRq
rQpjNkGMOxuFRCtwItplyjZDz+b06xfSia+u495ahZrMyHOjcXw8jTnbKPY9hhuPjlZarqbMsABY
VQi8Q0lM9bYTNFk3RlhRlHuN4nxx/wsYL6awDOyf0EccYaKwLj+3UAUaMfsd11nPRXZq59TuN1mo
wc6mfBpxdKV+Ec93po1d32WeHgxckDfVS7PlZAdiRcmzS9zbEOzIwLxy0PQ2b6AX9erEponvC9At
0OxLG4TzuCxu3Re0ybkeDyej/FXepdwaHqLN5kvQkXW7klM6AzM/QbyVSbOL8Bdak5tzl58Uus5q
ituNSu1nu0FqX611ik4GNmwfN6v6GYn2lgoPDvpkNg1Tl6YI1FXTbK7NNh7uqfUA8eTqBS5kOLr6
gwQUiP75XY81vUxDWcGDJbolpAlIgzrgRXzyO/TUeuMNhDH9j1mwnq4yrl38YpCv8zX521M04E6j
nWp0eiKIxfbUuBNN+mQLuzt+UntQ8XZnXoCi8PBAaF1ir3aOm6PvdJD1ww1Yt8iEqkS6sAWAtuhR
DNBXemTiGHsxahz5YZTX7ccD/9kYfEXdSJM0z++9CbNtTaehRMJVo2q8PndkGlijJd6487QbTt3T
RTV6yp9kP47pnBnXRgZboPDJgbuNfUBf8WFMQvW4XyNwfXkrihYzbNTIdcMWfJ+Q2PLcsjB9Gxw/
LHy4W9+zYfGZyeTwQRyYamSYnJsU7hyTphPWsR56/MhXjm8drogYGPT8Lk2vQd+iYvIFm99eokIk
dEkp9sc/1A3jeP7MQkoCjqkoDIZFe4F5CrJ2LvJWAl5xqwlA/qxa6rwm8o9aPzGtf0wasHNbudp9
gtsQIb49U0SUnDxS4XBylGSSHfLC90flQpWQHDp7M1rwsYkcvDZ2x7qxrcQU9rlx93mvEmcRxYbP
vxMKInFP4uSz2NtfizPN6HOFQGEAMyaA96hzMW3uVT+V5Kf9VBz6UbjxBTcbZStGZE3v+OJqRHMM
9zIbn4rRm2RWcF/xC1eOvFt2ZzGQ3FS5xy1fLhXbRIckop7zgY2MbT1JzZ7YuNPyFofEdQx9ipR/
P6ncoZGFB+HxTQd4Jh8KATCBjtGw0FyJ4UkUDf2VB0TZvpmF6nyxaLmWqta0ufB0r4xG3yqgliMq
F/hioMUjXRkkV1Qe/ZVIEm9jEOUJFbwsaVzshm07A7a6C0AWPZ5aowoU5WUklt6OLfGC+C+VLJgO
Fn24Gd5fi9Vn63Y1rb8BH3h2TM+AsTpRhCW1mfdzPTiNaOwxo9MAV3mab/0VRnNlTVZjtIKtNpi7
lQ290IUQGptWFr6xieoS8wDv2THwPULNnCa/UyzHcQs5wJgd9JR57fRAluw/ihH3piluYlW80Cxp
vpY2pvuyJN+JLo4uRWIPcv7Q0e/EAnmXmGbKEy/SX+GaJtZzddJUaccUSr5BcbCRjfh7vyvXC8rs
HjHENi9IcSYXbYj56c247IAK8ZaCeeZeck4HRqTjexWlehTce/Bxi4kEAMA8mE6srC6rxJJljU9P
jSzofW/xHTgYoSd62BUsxK3hs4l1zKzpGCDb4B76jXy63Ok5AcGU/17lzXzG1RCP0yOM3dAsBMPm
QwcUIEd4k0j1b9dUMfien4jISu8H/1R4z2s6LUb3oxC7FTjzdC/NUZr5PJDGemyFuR8jWr8TcWNQ
XrDwth06EMJiDtZrEd5x1BOrXtiJv1YoMCaHMB9UAlksQXqRGaI5AEkhwCqy17YIt80yFqedDHqD
l3Ckabr+Thgpr8kNfgafChsq1IleTHCYehFfZInPxsNsdT/papi49L/jrif7Pc4tcgN77CL/CcUP
pYNBBqtCKB/pUKm8hSRHAXlRNsH3XUSb+an5cA7DyV27qHi0ynJJ4wYTpQXJztDhE19V3UbGGI6t
pNVJuiH8vVTzhliexeRVeax+NBn6sZ5NJCEXQShhRzfVHhdYzmlOVDskdw3CIWsmypekDM05neJQ
lOxu7cF7V5IvJ8AYevjeB4MIaolHGJnqxXe0rL0Pql5O+ndMJakNJYi31s3l0JNyHF94xe3jBQ7W
2S5X75+lyqF+HuIL9GTsmIihjw7/Y0dlidMRpzH1AK8GpxbILrBIcmHcHeiJc8MZVF21aFjWkghk
iUzuMEd7l0vxAbolqeAJCuMdgP/QxlvvtBeOlzQgZpFkxX/OPrY0vNej7056i5J1R1BtDfrqL+IK
KPunZngwW76A8MlDD9hhGAQ531uW+8lUAnuhuqLefD7QvHb934IpjKsELfkMHSopEezYnrGHO3ZB
kmdTVkC+/HVu1TJTsfbE0hwFKmimdvDZSjU86xb9GLj5T1UhVcbohOU5NWLqOXa2mIXXxZz8OUvw
PfEzjWLdh4UsZIYElpGYdamSk3cmSS4VAju5J28Dtv3EG4YwCsavULA7bfAh5LOfWCiic6ctpcN/
S9+jZ6v3yRckBx4zTD+JSNpOU0uYjJG4LQ1gXfWJ7Rwa/5xNQQUNfvBrcDM8DMTl2n58F/xdHJQR
0UJI7n2A0mqGSp4PISFAfNrQR/m9HxYCw4dcXxRySXrJBMCVZERqJIgM4RB9TMcs9b71aO2mQDTc
corU6qiG5c1MTlzeTAblu7ZCW6rDrq9yvtRB2ow7tFB119S24fClQLQu+2uLdWDaNRZjtbU0ATLz
W8zRL79O5MnmdbDtKLWRsRVUnVFdfm3n1v77dE8Q+wno9pgRJs6K9s7F5LyQpae2KvdmC4orAXn2
hUrNyiEoiaZXe54svlUMWc9RBR7+5kSu0AjcOordnnN8pqUyhbaSTBUPdOgf41FSCEBWz1+m1wid
anHbCSqimIcSwlUXdXPBLt0fB+iHV+lSe/wODLUqC3ichHEXxfw7dxXEm48xTmamXi3ZUz9qxsK6
h494Mw+eMvme2KqTAN7u/34Kk0Soec+9Zdrs8WYN8gIQ9BvzP2XM1wW27J1XpNR+5gQCpWQKBsq0
e31w56Xvkn2L7+l6bcaEoRQDBtVd/GOv2SKiAW6TZu/62gxkMXz6xwR4rQoyQV/hcBKI9F/5OlzQ
hm0/stT7UJQZauiNuaJBubbBrSPeXRZ5Be+WAZAqcxlQkZ7UDw8N99nc6EArAjVaa/9OCncMooyv
MLQuCTwB/PcUzOgSVaX7VlqlhcF8u54Zt/eHXuu4RdWaMn18hJYqzO4HAGrc98zHfLsp3hhF5K/o
8nMnDOvMCaxmB8fXyRIWdAoBtaAjjF5/KWwSDcJUKFQv9hbhrgVETa9cE7g8clPapHC0aB7Wweuw
yMv5G0lhXuByZXue2crsJQB/HbcJPlVNB31d4XUJn9nanO4wQMIFVWp9gMFsxFnEqtPSYZxJiZAL
a/4l6j6lEIPaXwThBjRLaA89jg6iponkAyXUeVXkmW2C45FsTtD8P5UmCx42cKUH6Qh+6Yq8FAj/
g6tWLfHH+onHWW+RhMZEBQmCe9H0g0J4BbiRrMVMsoa9My7A0zJCcPkEkJhFMWxsG6ZsvGcYhA37
O9bhQaFQaPyLrN9NMJBZVj8LCdCDpQwOVQgqk3gNyR7LUB8RcUV43Wu7R7tuSdsnEjEVrXNBptB6
3zhj6wnDh+U4kWNGLFjvkgQf/ak6c8KRk36QjGBi/lU+ULSdNiVGEMrTgW9DnMUtnf8QC/nkbbxM
U5xh72AYR04UjSxdJ+GS3uj5pIzdEWy0DksOLXTCc+QS7cxTOh52X7//ZpmdwLRgSyc8Ew4O/R3x
YtfZBGZn6cod51lL3JK37ugUypoVU3gIHPIWE5ZLBbD9ZCkvo5FF2r/8sILbHMsv7eYjUdXBSdR4
zgKlxCfZr7JPW2EgiXpou0WS1xxQxddwDpIs5159vGbTPl4k1srmrx5t1hUJ7Q6k30j+s3DGnSDP
lN3ZzgDI8dx+/DwEpLjhsK9EqJUyHM9co3zmta3DITL6mc4ten4A6s2nvy63qfftjrq7EkAu8xhJ
iKMzMBEOj7+RA8vUcHPr1dTVM6TSlIIm6bOS4O7PgqRryKInATzjgA20VxZj1U+fgkSe2u4LqorD
uTakAVbGbjOc27R5pBzRP+AQ90Gs+8ZzeOvqeSt5Kv1q9XVTof/FZFlGa/M/SANPGxOpGzOmPuAg
5U87ksiHRI6oVLmJX9ZbmesX87NVL0Q6P01wXi3+gFHWXfEnqmPqXeuhP/QHKPINS+mT8sSxYxyx
c64R5W1OJcxegWT4SjG3hEWrGJ/O43SxPGwCJiRGZDwtxhNfu5AQ7oFROAVTdygp1Urg5ACMoUZL
ssq8crk1oZahsqmd0l7KA5nlD9qMT/B+uK87crIu1JPJQLW0JVTgBVHW8gie8ksfZZA41olEo7aR
dTnlG44XhnZdv6xIKwk7AoClDAjJtBJIW24A2tLE/DGESKtoqcnBJo8v3Kyoi9kR202f8e0LD6Vi
HLrBGJWV+MviAAdZLve1gUd7LtJ5SGXsPolmtI6bwAH3XJmBXmNM+878noyHK1X636JINHF9pjlR
Yg0mw/TFXU2ZCUiuWB8m9L5XlLMVEytPko9fBkQgXRq2FFl5lmNDSYMDK71xs8pZn1v+yiv9dHp8
Sys/G7onikcYq28KszZu31Ojn41XUHC/6ESP1fv/d3hPya5am9tqFpspMrSSYWShuA2rIwpQ6eXq
Vzq09NDjTyKP7yid1w0Hh5AjD7Exm5uCeE+iKulgDzgDdhaae6/ARFxTHLE93tHI0xE51uAaM2hu
LB2ZTgPO1ZLCrrn4SCraR0YsKBDUQeCYb2y2RN2tFF8ZpDIcCDdpF7P3Sy5cp3XNmJC9/x4ymDPt
1yVFrZDCynQSTfmTzSP9Z+OXfiXShWKlIXu7LIGqV4wB53DQA+aPvp/5H8r4etYQceTzF81MA3fC
MnrChEnvOMLEFDY4XelL0qznf7FCQ1CIWKcA5m25qdxJXrlqTvszy3BVRldzGhOH8wjEb66HnHsg
g7aKQqT3W+PBxfZ4efduL+8Ky7tsrMptfMKqMedNrcKTp+X662FObvneGpClzs6WX+oV3v5sfqMr
e6o5CyRMiPEhGaNOmiAVgiDQzjy3N23VcHv50s/nnpt+ub3bqk9HmNXn8TokJuQKq2Xo0VJKGexz
rstH6jSx/uv8JYCXkMZOaxyW/q8YnfL57ogsTsxQOy3p6Ed42wJkXnf2LHJOvgtGIdpgk02Umg9D
f5yBftSw+XXKRvsEDnenHm3+V1kXp7p/6f7ln8QNsT/lSZvUpPRfs7+yu5kUWnlMVwPfZDo92nr8
mCglEhwsb6EjBTHdMfXz8i9AQkq2kbg54mbQSISgbP77z+1a6WBhlQfgH8vSr0sESfTv57MeS/Jz
Xg/gbgK35EMdYHudT0iaj1/EnZpnWYOEr1RaVUK2UbhPr2g7IduTb/bRxxJJSP7qPpYChzXU0daK
vYVeUXWipsrA3nQN1iXz5fzOkPBAXwu7TExzBA0HN222jV3CvaR3yJallJktFlS7zjy9snUJmeEQ
qFge7Fp2nq2kVbI0u29tpsGP/qUczzRCRfB4qvl+jYwcuFyiPb4+81qkkxCv4I7JIBBkeqrYEIkW
LSGE15dU/Nc1BZL/ioP0Uj8w8wUNW7tjx0Hxcc/bnExOqqhXGx3eBw9rgWflAeVeVwXrVLNfzU8v
Di96hTEOfF1dhALbdvkb9kdsV/ppXGmupOFrKfTOBB9QLZ2SAzUhz7phIvH+qruC7Y3C9T+wempI
wsuVhfqyXsIogFs1D/EziqfF3aT+NBrMPoCW4JleBUNxJ2WJS3jZ2HoSbD82ra5V1kQb0+os3bWf
sZx/iAKF4ofL0o4mj4dKm1RTWM+5Z+0KZagkWD7eHjqy4HHwCzpTkCVM1Hg8nnuRHm+nSMGnDdVr
NsjqRqDp482q/bquFAQ27piNgEEdY7NZrvsdPqLKt2Sg9jG6Xs13dKT0AhFvZ4QjNXv+j1FcDc/6
nJEIgg5xcKAgAI98G862q8/G4m20THyi5LKpvDh9vbuUAZl8fcNImAaP+MFdjA2+5A4Y+2+2/gHo
2i4A1fhdy5DMOFf53YaP1Rmezd367zJM6r2LUONj+LOiavwoCMtBqCAlw4/UZqcgWeRiMMSKj0jY
SjSGemE5/JsIa+Et5N0NRjX+7HXxdETEv7vM3AafHznKf2bX3UYAy6VlMg3G3LAoFF2sfK8zONwC
pw5h3iiT8Niwqdmes9Se/rv1Q+OovYrcV3VNzCWxgfVoQhanCKF8dQltrl+h65WyxbZwcPF2EP+b
X6y+glxEQAr+Ua8Aokw0uLaI6YTaXnXB4lUD8ZHw8zV+dEjEs8QPd1L0q/l25EEmcUun2PT1Eb7J
G8uuqsjZ51m2JMeslHdFZ5VOZ2qw19Bn8eEoFMcmTWqmO3RXVsMb0002hhTe6T3q20icTWTqR148
RKGjWflaTfkRjGrci4FvGGRCdhLC6YJ6kGMjPFLbIMLXfWiklWb06fqQfmdHYMJRkowgVsYW65QW
G8yIdJFHV8oONdzUuA4l4mP28mHEP2SicgSfLGm1AUIl3Zf1awcIBzWt77mGa9bCfR/6McLd4ys9
2WVjuE6/HtRUfj1b7MmffFLAXhXetXfBqOHrnH6lUE2YHMfsLBpsBWwGmbqORXWDVsuxqoKz7GMA
AUeYxbDL07DYp5Mjw5MHPdTxAYzVOiaVMg63uGd9e8I/1P/fq//BjKrRaC47Fk4SKm1y8iICGbTl
RjXwlUIEH8l4vU3YnOai7L9UMBFnyeEnf65falnTOMTcJHCV6A3ZFLIQ8ybqDAZukXh3NxiqMDnw
/MGNcxLSu59/Jp4ck+hpkvEgHvn/vJrGS3BxlSrluxYWzT6i9UQG6PLNSEDCI4P+wxHLQrDKpC4M
N3QkLdl0i9qYe+Wt0cM2MYqCytRR2XHvt1ftF4zsCbYa+BltFdhIX0z/lGWqusoFNLONoqinBQEC
TJhrXN+EXyghwKNJNMsHJutWLMq/z/xeEabaV+GvODCkBHzZFNiitp6IR5yg/w+uBbxbBW4ELbNG
obI3QC7GQcSWSlcomsI3rw+ViSOLBatnqm+M9+O75UcG9pTTQEFRY7/HdVfq6FnT8RiRBa4QAlSk
TFDQ/E3otOVcM9GFd44A1oYrKLeN+ebp6cUhZfiKFw7zWF3dfgbZGwLtys04frtARSQSO7oZdYcG
K8NL+ZqI61abMvYPaKkriILUyU8KVwg/b+d4znnAekImS+cMk6Im4WojsEFccyPqrELxdsXEjzKB
9XW2jqUGc6/Y3UGw8qjW7xILlYmFUA/Qprr7yzFla+xxgkjrXDY9dtlTMe8Nenvxd50uVTHq0hFL
y8964/S0VPf8y9rlrJsM1rdB/FOCHdsq2Mi4zT0ZvTvUzfoqPcx2Vr4p4GZDeo0OoOzUMbskWnwC
yiCwMPd0wqqd2gJmpk6ir8hSqaVQtDRifdQIeqmbxlJVueSEFCL+YkBPmkCw/v2xoeJHZiaMUYzP
jG3xR5w2ZRXQyYtr54YKxuYZGsw9QFka4fMhL3VfrIjuBiaWr0e1xAc47rx/kWToeWIOn5ymzmWZ
E2sAcXtwXPdP5HKO/h9jG+YduPwm5awy9nebITxSSKiFhQvqjjsTz+r8eumkGQzvX+lS/vS6bEmI
F5oHJADxP16RQYsB/rRxwaJl746+uNCNsmwXYtKVjfb/7sP7sd4SPVtPXBtN/RoT4nj1qqEd4pdF
2k++V3e5u2rQLXOKkgl/+Sg197ify0+YAdKiGszbKhfLWMqynPFyzOolVG+6iK2tZ9i/YvtK1zw+
7vth3VnlFLUeE1OmisYSBl2g7xbrnhIxOyxU48vsW0f0sALjCG94znLJlYkE69lu6GxIJ/Bi1oxK
m4S5GyQlFcU+VHN8PPCQ+6yAHLylaQwNZ++zpEOiiFiHIKNOGxcA6VE39cUTcm08eutizFKCx/9p
Gj4pi/F/UKh4g66FEjyLSAL5Y4+GedzZ6b1hwhNmwne6U7b9eglCeKWmxourOHrGUFf0dGzBhBlD
VpqgeESjXDtM3nDezzmA2u1BynKHlt5KDxZOR4fa0/DYJ2Jc2kDIVjQFVfe6fpwUv8Ff2ulTcAi1
FFyBsDlfLDOn73L9FUdutKixjUm16gzhx8BO0s1E5iLEwZo6c6Y1bUzRZqWAPl/V7ZnIlwu2AdZG
xmEr5GhgU3YMh6OeB4w2ZRZ2URpFvQe783AYQewXeqqmT0GbnQpqAT2YA69F81ee//F8BBva46Xn
Lp+Luer4d6j6QiWJKFDObc/bD3RjDRRkwgB7uEHBBi3zI5zdWz11pgiqn5FEQJYwTMreFUUOHZYi
vTLLPjlCopX5ODVUVBYSAS4fu8uXlZjrFMijp2njSHOdLt/+IQwScNfD4JKNGXm5gPshrdEJvfB6
Hpbm7VrB/tLB7QmnHLv3udtm/MB9AyMFLXp66Q7cLYeDxvws2LoCCT9NcuDsTizVhMGgBT1EGzQi
0oLtBTlYxzH292svTxfwl9sVohKQIlCB4vlGK4cahQQnokDuswWqjA0tnBUUWsqlRicLab8OYp9C
UcrA7RntvJxXtE8M/3oCFmjiofQtatVmzUi84AefUlIaZ1Tti9FAcZgkDP1e/rVyctyzFjB/1vS0
fwNDpp0lKm4dZ3oCmZxI89hNGvtGOT3f6U/MqNLDArgsFFdvRRBb1hBZjIxz6rsm/fQcVI+DBanf
Ar+BSSBHttx/XPvldjLsDHVjIuQDqL2YAWc3Mj2wjaiuAqKrVBWmt7B0cAnNq5wyi6FKc+l6k5cx
nG28SKrmmMZv+mL+XovvYOjNSgtMpL10xjfIaPjkMWJybpA+P43yj4bMsId2yKw+EbEV2hjgAWFU
A/uDkjzPN2Lca/5A/0Iqv0PTy6Y0/+ZTwu+ukHpR+YkzfGjaCTdZMlWKsI0eeqA88hekzSt9kAQD
Xv71ERwL5lozqz6pUlEy+9XkMW2barZtJ9+f5fxy7kCxC12WFPcD3s9KJg2TPe1ZSJ40K98PyQQ9
SLXA7PVKy+dk4WtXQDpqRyRp0ObdeNGTDurO4vd/Q2bsUlKtLbPw8MTdxByfLOo67Df0NrRd4L/a
LwdMJYwDk5A50V5mIcXgyPh3FA90QwBwkjvaF8tZinUhlx8DHikvIj8+ydNiK45IXTXXtWX8QiAm
Q0/x6O5fdXBmnyhBoHua1yKxAdpgLWqZOXBN/vIFEdniVz3zTM3UoMgq8Esp4yqB5e9bowmoOpM1
vPCv0ovpL785UZgKT/DpgVZsKOt2ejuMbFSP1w4SAJzb7epo0/3v/q8RpZkWezi4tzMoYP7pOmjJ
oqoBppCEpY4YEzZm5PxTezIs/iCyJurH7unsinVueK9e/6NESU6w8bzbMIf7e1ePZiIkY99/dq0n
4Oh4aFtDopfe8XbK7IqajtkJhSpfUMzVPEZdL0NUGXkUnZjjoU1B3HAuVvXG4dsG7D9lxLkZwQei
bTBn4WSOtp6XD+xT6rL6ww/K7xCZzPfbGqlK3sNdjMZQLKLNy+EjEFAdVtXnOlwrhqxlmVu09ZRD
BYhfcH5XZCR9WuiqmBSPcMsB9kmamonLZxQceDfjMW+pwBFNIs8KIhpcJbKQqNM7U5/4+Kt2vZH4
qgYLJey95f4e6qZGxWY1ghjOVyQnx8YWgEeeEzKBcFKe4AUVdYppeSj3FRrpVZp4Ol2IxIBMqw26
Ch7ef5ZWn+9uC5G7dBN3nSLs6EHtLxzbK8rnMej21m+z5P+S66yk8sAOgKdYP5W6Xk8W91dqqd63
Hfz7J0fKQWQQ9i7y9i16Urrt1TIkT1qndbPZyZfKGXCtoG1uY6I6xYfRrmqfUroDF5KYI4OF4eCO
l50Ri9ClccehJS6gZ2vBKIJBsXOIycLVRAtNjIm/9Nu1oQsbqM+0Kf1thiwUCay+zU9u+Sa68Hbf
iQDu9Fh+HgTWm/QmZOw8I8BAmGJiUMuLxiLk6v1Jgu4lykinpJgMTOPjzwL48C0jfsYvLZv27dmb
gyIXIZhuDAH9ZuZM8EHxPkBgSXbib0slcD/SYEoOdraroATTFd6RptmrD0KhrdUlJCewNfpMeWmX
8MneSd9x7MdVRzd79OAT6RtQUn9pU21WRCV1vLgQH1cYfQ4wYctmdMRiBo7nhLea2bRfPji2RKU4
15fkTC3rlwfalxoYAv6NwQiqMgNp6PaXN5WKGHDKPPGNZMhnVkT4t4qYVOmGSBWH4s8CF1t8eh9L
k7EhY6TG7k3vMI2b//TBtm8mtwOW4P4Fhfcd2Fcr9iApO48JYCN2x1X8FwyMzEYmrcXbMdc3QhX6
y0ibbbsNlJIwcX6II8gDGxAbPBjSCwrP5Y7BCZ7haEmFisIJ3vfcFRA33bVA2cAtjmviYsDv05ez
wJ4yKGWguW4d/t3iBDDpn90O6seFgahPMHqKAwSECtnDJbGijAAfM8S3meoNUwyDRmDqKPaYIJ8v
u+aMjJIdyq1anm11WubfsOQg8/bDjS9TqThVpJoCpbQLyPpTuvopgHaEsXwDfS03yOWjbQHzf8w4
6v5/9HTocvbIDETt/4Trh8ktW61/+9qKssYBjFZzTrkPmKVVPQp39n43gReeqVbqqGSS6nNdS+BF
OzZRRFbbzhry7nTsHXizkQSbMnxR5j6pvkCcVjaRu0mxjN7rX7BQF60LiH1dbpltexCbdVZX1rvy
CBlWD3xh6GHfL36TZCFGEbJkC/JzUyZ8xVN+LUkT02Q4nas6vcy3I1cIsj2FnpHzXbipDSeE+/xi
x/M+Fqt4+CjbMM7SGCJnu1071t+CnbWG5RpIWh1IRKF7gJa1k8qcZAYfsRPmGJsPiaLVUnTTeWfF
qXFn8+dyO1zr6MMt43+2EumN4uyF7VnJT0pML4O8DcV7nYPnOpToLfQzL4I+QvKdD0WVWVyFXsuN
+68+6B2N1Vvm7xf1XWzQ6w4tD3Oz/7WuzEjV0Y8lKbhfRAk9OgeZl/kah3UCbxpkNsvF/C5kZmmk
TBM+X4UCg/4N4lPtVOWpNcDa3VWXbM9Q/GqxhSQqxqZCTvDIb2kkyXpRoReRL9Tv09J1qqoZyCnB
qEk522qqV2YJ32z4SOkNJIVtAQ04ty5STPQ5sI7gC8qEAtfJpx2XFL6HZjwFI7VhgTM/+mh0D/HX
ByMF6mzNFSTtaw56b3/FOwWCDv9V0LQ37pAbU6ukKCdueZdVluGNntJatno72IR6rG1MVRQiT4bK
sfXqnCSQ1exextGa+dLXjiv7H4+F0atdzndaphYcjIhZ5VhDuJagAUEs3ddYZrF4QiXE/omYlrTZ
NQf0yU2rA09CKs3uLrFUjFCLqNZDjbzLQNdjt67PIHCXpb9IqOVsnPqbVm9/bSMPDqsBv+xr4UN7
vWtZQK33TOFJ3AeTw0O5iFJLxLetmpRupI+iZuwJvf6h6epA5Y3hqj6SgTRVRo6I10Y9VA1BbOg7
P0AzDV/ZoYe0YJiUtbrQMYx8E2nx9HHl7/x0n99ag+Lf7ATuuEjyhGLsd/JrVaGfPLX+2FgKZxTx
6iSPdrXOkphqJwbHoiLNTeg+yu+oxVPWPx61p44oXbgkqEeCSCAowmgTJyfnlqOYeSt8ZJYvcKvr
fHAfcX1sIwAE4UuZkb3nLlVfzxHv+KjL/wX5SJF7VEpm5TcPUNEE3d9PQsHQu9q2z3eMBFog9lpL
S3phTvw3fqH3SpDWwF1kGrXjwfng9gTcG2nKdbmxSQ5jDj1y4mgQM0USJeciQPLo1OzzHX+/d5O1
A6i10PLkZ+DdCyDn9zwMjS4z1Zur106DcR9KKr6ru4+4Zp0AX+OZ9OWPn2un+2XWWYzwSCgdBG6L
dBUNyWZBWemv9Q4Hs9V+lqs5xxqrMde+q0NyGudtq59bUViXdtnVO/3U4AFKhivpAb31u+RyecYt
Ac+eiUH70pUomvmLrgz41Ilss7E8AzNN9yV6QnSTK7sfmV/1s519hSO/LuCWILOmBUS7Q51w2B7A
13uAc4x1pw67EzpBI8yUpKyTRdLWsajQmVnGc9sEleTBS+Zi+yyD82EP9WNnamIJQeKdvfNjEhp+
EkWh1UGhdPOx+HT2p98URTnar1apcIZFEBfxW83JBGnoU36DOOhnqlnS8G358YAhRAhmsQUvqPV1
8cOZDglHNDP8qXG64MBKsY+ztXnZnKoRvd/KLlpmBXOhSbMFBpZRbhaT/D8L+2tsXzYeMvTdJPFx
0uLF8Q8TE+yW0yKKh9ySqq9XgSL7tf1FT8Fw6vCBt5D5Grf1t0ngkDxK3UklcV2X7mba8+8uhQun
G49jqYzSJcIeJT6P9FMoNAnl+IwI96E1bFSewMH5RxofdyRPmhdE+zh8dBVKtpuOuXnoihv65FU0
ZmNQkgjI9lZUqjlkmhp5P+4b04jpWuNzduSEijHsMa/cqNy8zFlA/Ye7hCV7Z1BP+RTC3AZ3qTuz
P1SE74g6/YdBc1z3Lj2foGYk+2q2DN1jVnr6VEjYYOvqSLI6kdys8JaQ28A2F3vL/wVw/Vo7B1kQ
tNT601n4XCvzRCuHkQedp6bcvoyLMX/xkPiVcoTH1cxyNAp3HF/FDdIHiOIAE4EssomBj0l1Fl/f
F4qo1YKAMfNdGgD3VJ7bT38/UolZKfMqH1DixaQ/QLW75wWZXNMuwrk6JQW37dozCAOpxNWiavgo
uOAWe2SeLV0CQwyVljSRpxNA2hLKYhu/vWmuF94D7DEEbr1ocHu4Nl+uGtpQ50kT34JKzgvw/CKr
z2LHiaFAD6Szaxe8jpQjDvqDqrnYC0k49YyTWk0tqQ8I/VAaoZfvsSrT/XbqD0EFFuDpQLR9tkOG
pahXjRounoEF6g2jM+lVqJgaJCqhjznQsSYXXcQtZvYZJd7/13v/2qci+SRe3VNJV/YqDbFqs2es
95W/GyncZlAOQVLUQbBdUGhXtM7p2z9eu3C0SqoptiJT9Qzd/OoVLUm5lMHZVNzmWknVtfZaIZZC
Nep1k3JwjOGic3dCnMfAwUuFl4uNg5GbEzhn8NzMU3AYUlC4JmTIKCi8jp6ScJNL8HTRrCAOK7aV
UBrDrUZ8+SDydk+/btpasJ7C3T3FkIsZgJG4RYsGfnuK7L/KjjHEKfOlaMxd6zjCw9t/JQsKjKtr
bI4IjpbWoqooK3EJ2hwklrMrVDne2SL9k4edhDm0ARTCRBKeBo09FODayx7FZwMA5yyH+fqGzcqV
wkI3gj0q1UPq6OB1sKkE6nmYM07J5HN+zm4irr8Of/sin4nXFZ+99I6VLnG0qUcsQJ1NzzWOuRZl
jnnHggqSD2nQPBHnQqa/BWL9DFsJr8xNG+tm3q2+JRFzcHP7unV/wkhtJnO/bIhbhg+3/C01jxxD
s70IpMBkWVGSGlHGi7ToxMgoDB7PCL1Mo07e6LInugT/q2UEC4nLm4VBftfu/ahCssXjAzVKzFYK
h9gWAKvhOY4ZYBg3py6I32Y/+jraIhzzsYgb+xzdQrPLp6Tkf7guUFljvPGeWXRdlRYI9ScxeJ1B
eCV86/D96KZJWPT7zMP8vxS+C4a9hVz/prEfrZTCNXMIK8EngYy5/h8cQEUExMm7//4xdRlm3FW6
j+tZC5OBXEshpZ38Ph7U3jJBKxKbv5hwi2Z8WHM/Z56bzz7KgXgsNq5xHv+hNK9o/BOZ3DLAMmmM
+rNal//eCmBMyTrlJYyz0ZIMFvB65bicodNWfhNYCQnbMPuRIA3JbX/9bKQY0G9QqmLaYKX7hviy
6SukFsynPCial/ETBn+5gQrFcdzuzHigu6xC/VErFBWDRTCI0K+nzgIJrBEhnd12+rNJ/pXvHTJv
o2yzY5yu2KxouHQaAA9b2i3TDcFrgfi3xEyhGufxf8WEPPuu5ujPPc+jNkFbweMkSBzagZMTloEw
xkQWoJEks/BaNB+W/aUxf2RJAEbYG/Jjh40dDQ5h+CQG3KTM2APovczrQxUothWGsu8nOvLb6aTb
K35ulX6ktX9sMYEl3qvxVQ4cUvE9g2aVG3zQ7UoPwlBaan5QQox69n2xmTj+pMUCm9jCb2NueSny
nlk6bCS0vM7xhBp4ekMIhxffeOvMQoA+FnMiUJNqKXJVzz1RdkswCi5q8jvfZrLmiJBk20TwpCXL
Hk52/efzIj8lZihAq1iK5k0c6SO80EN5waNlC3/9jbQhxDM4+6zlS1EsDjz0SQizHsdTqcSefpUE
7XM0e+n0lHCTwKYujMFY4yBaSitvyc26FPda9U+ft1kV+8rlqmrwKz5XMQWKvqFhla6evt6STiw/
cDlKQfVzi53PShA/J9cUxyJFpvb/HsDFSO15ZTfbjbWFWuL8CM4+nqexdp6aYPadVIfTClk3CYHK
e3Al055pfPqg3g3zsn5vx8c5aZZbGM3xz6rNa3oaTYjE/LW2feO3qGrVSumZjLQtS/Y4TKeICszc
VD5hZJeyBt8jVUi+Ik1lX27TVSr1BPcLzwIr834kuTFtAsk4DSWZ4Y30JhOxPfncqm2G2l8cIlw8
tl//Pi841aIiHjQ3Nt4HDZx2yX0PX6ZnHz4qc9+XF3usofOJZCFqUA0vIpmCjvuvgIOMq20VJxGh
lkLmzeUCIuPDEfUtxnz9HGdKmhd6ppc2U23gA3WmkQ3IXn9NTkIEFg+Odj1EggBDi+3YberUCYUI
6cI4C9FZAwtM3DKEOvjoAl/3Dyc8nYa/qt0ElbArkML+2KCh14MIFsojdVuLZ9gEeBqbyNCsRwo+
2C0IZfhvorxWTMe+/fjg6IAOiZQQl6qCx3l2axOhNYRHzG8Bu+vOGjISHWi079PHdyzEXz1YgphW
HyY74egx59u494C7TvHdm/WrH16FU4HrXCeSSTPZpe3v6qngh2cIRZvIlV5LCiYqq4+jF4EbMgms
NEuki+Wp/oi7YGzgjGt0XsRRYjpDpZwbD+LLP1izYskTgI/gJW2F+JngPId5soAEuz/lM8S/uMKA
AMzhSr83flgTYNImrPsZY5XSB8TfFcIleK8oq9PZ/4/HZfDpwzZi+s89wFSGbnH29zLp3tnT6qk4
GRGEOfedxUzryO8oUp+PCqzgQwh8H9HzX7uVWjSblrawdKRQ8IN+wBZCCqr+Buxco6YNpHhXkprd
WdPow1e5en//jB4dnIFwz7Ukr+6tbCdkiqXTKy9hzOqIXeaE4SiLObeDPeKgfTHZfYGDngQ1CA4Z
W3KTEDQxbTq+libcca8D/Pmqc+h5tXC/ouedDawe4E7IZ6xm0nR1lXbmSQP2YnIzgFO4F3o5N5zc
9jg1dV64Y+EBzzEVyyXPyG/uCGkGMFGBBx5qeiGVkPBlFAAPvMNDLtGbwunPfydrbMhPeNr7aD8U
Bija+S9ELLu19UfOaBpT4QlUX0Zhd6lBovKgGtMSQsylHg0iS89Axpb2XtO1Mb63Jrzh/v8+xxl3
yIVKoP9ILgCYXNs5eOSFim3T83XqrmMsutRpfS+xeDp4bgt5n//zaWWOvpxnfs9mg40wwqx8bcfu
lVw3nxN9HLADcaz+oSLVZ3PhdN1iVGUGR4PsA0y1SZO4oY/GLCf9LClpGL+ocdExIObZ99jkDwKq
vF0LyjQdTBgVVZyjvhtP/N6+LoPfYgz6NrZShACHbOK8+LSrvEiZ0JL8DDIW4SLb/K6HaVPKaENl
2etrKylIX3yQVX0RbBhruOMLDLmGMLkAxgd7G5HP9F2ZB1L1DowSbLSpqqQy1MdmeqnMT6qhAqSa
9WSNe1Y9+PUn1EUyOkHHyZLMqDL0TxcpHsKVenUDBj7p7vAGE7EX6H4MYbDibnO0bK+ttkH3Zxml
XSblUCtlFB68QPuuwFjhVhtZOjqmv0p0GwiKaqEkDnedxF7w7/sngewEq4ieCpjGOsUpKdCm4r8g
7hCPIDH+Wb86+QQC1syHRBp4FhpYKExXFG9kVgiXo+1LxT42+rMns736y263FiMlST4fudQ7N+nl
SlGkkk1/6zlryEsKDY9W0lHPL7cYYChlRULyo+vIJSjH94Q7ekeNTvAYxYrNTz7dOVb25pcBiyy9
wGHGSWf0ZoVnwECUUd0qBysnYAcWeoe9Hr+xQenHb1zKSHVJfAZDTKQlHSxyfF5S9U+3JhX7jRrA
iIm1uoDjUGOcXLFfaAIaD63rbAPV0G9X5oftRZd4Iw00UZ7TSN/LQ5aRG9vJ2z0MFLSgIKG90xzJ
nRic0Hw6qk//m/qz0vWywmI/CXrIrLzNYgdCIs10gQHFwlvADLxguMJJEiRjSMcXa6n6TJ3VBycN
GH1Z20Sw6n+9WFCmWSUDmpCrrPq02QWL9LVFQgPMaq4J+EmbAwOVWOJC+5AQ0G8EkON6GWhpt+oW
5uObdLqj3XB7kiyJp++FE9/cEvy96xtXbQ2b7OQpS4C53JjOsh/OuMzRVa2FBXtnbNGDl2nTQi6D
aDW5KQw/KK1fd9i0bHLN/C47BMoclu7k7Teg0pbHWVFiPB9p5Aij6gwk0GuEJ2Sx7On0Q9bOkiAa
qUK1E3vloqWAhjH3mTaUt9f2tRQ9m37gYjlKxE0kyeB0sNVjjcsseXK5NMpDnMVHpXaeOmyPW097
U/2bn/ZRjKkrBBAty2C4fHAshTWdBIEMI592iDxkfRqOqKE1s5Tw9wpbE8hpaAbRhw1FWwpB7kth
o+35iJE5oqmNoJqLLnGhGueK5YueWA8VE7H0CKOs0kqUJb8Siv/LkUvvMffxmAux2o4etcXqJ7HT
sgEaZj9JjgYsH89ILu57C3oklIvkJS5EIpaKwM/bIVCXFg0t9xDKkfPtAWqX/GuRBFTQefaxs6cU
x6j+6AbW0Z4HvsA2XGr7CoYHVOPWhgAOsGCEPZU1Qk35aG21PNWa9iEbNgehMlLF+8ZKsCouHO1N
2rM8kFW90q3Tn/RoG5wHpaj42Dr1+8B1akG9O0EuljJDlNk+gFddUz0WjT4ob5qu4E+yhwwk0djE
pEF1wt7aO7o9gRJNYYx5dCUeD6TlJyQ5jX04oWkHJeAebo9j6qwb2n4cbP6XNO5ey0YEEOXs2ACq
9TGbzVAwyhDHVNDZSBkcJYyVfjImBvBAbOPQM+2w2X4KccclQIlCm4Gqe7heiOZX7OxwgH4PKbhm
7XEyta3uQA+Hs+EmhVRPRAv2EdqusujgRgqw2eGLKTqB3ipFrpOIZO1//L2EW6khExc48Z9ANS1P
JAFnmG5HJDgajUK2SS8r+F4rckHiGGHCitCQNfrPVXIrr5ZxRqkdSrLh2Em4z5rSG7PSxsyL5AoI
D/B3Hf413fReQuy0HriQSbAcsmmw2l2c2hAikXLUH5O+huzfXfuuWhWP5xTYkqUM3HQwE/kuJuiO
A5DmtHSw4leGRWV1eN5CnMxpe/9CDkv2vgfHmi1xhPRjFi1gLln/gOkRiS4QNNh8o8WlU7BCh4Pt
iPZca7tqRmpP/9O67pWtKcTuEgLTA2qwAvfgDgaugbIB/aYPWl5WYmijmE+AHgXxjsiEH+FkZ0Qw
G3I4a502bmIt5fEHAMwnKYNSonEQQCzaQtkbxisS5HE1IG5G2K5wT+l0qWeBLOQPdBM3gzS36L6Q
kSwzyOss5LBnwo43QOVJXGru1VBlN5OnKHWnpGR6bgkOohHWS7xAI60zuGSc+LabdgGIxdbbNM2+
84H7RPWSPDCCjC32TKra2iP2WsrK92FlzH2K8YtxKc+BJtIHJ1DQaUcLBMP1zocj/vB++ODFpWBz
5gh5uhlmlqdmUHoZLko7/3u+GNcCpAYz3QK4gW/W6V42JAUtEBkjEpZqw5I51epYbgA6yfQtiG+X
INJM2lfMBB7j75cwipofr3h8QbDkvBXUoezfgQsZdLleC3ClD0/YT0VnGgCrZADPGrOuqpmTjhKk
WowQWiUQvxDYeM18MkKCR/WSm/1HbIsZNo50KQORQRxlqdSPNCnCytUu3ZWxv3hFCQKTImr8koPN
48ZH75r41NRo9giI+t4lflW/+x/H0g8Q2aOLsq2wlhUR0VzWOMM9sZWBJcrDDS6Va5kjGA9if0GZ
M1U4PEDQFhDUDKL99KOGMWN2b0bX8tNQhGkSNB7KlCdccBnCbMvp8fW/WJNFs7tGkhhYasdvLDb2
uaZq9m3Ncg5zXFdNqXdQb072hmvz4s7xAXte/VwQE42Gy8/3JVjEEY/actHcEoM/8cRyjCsPSP8G
cGP/AeEvkGZP4tkcqdVwIZT8SUJNIRduwJej6Iz7hL8T+n7yrFbBYWppwwiiBSsbfxPL2iu5Eeio
sf7lOVXc1IdAQmDEG/Hw7Sy5mxbJhadHJRQJVIRRevj4bjZ8D8MQKTwLrRlUspj+oieFkdYCcVjT
ZBIlPyztPdKH4uQdtOCC0yiPEP6Z76COpxWM+8bLt6AcVIfoPwwTkLh1tLycerlywfyPbB2xuoql
c68Y1CzeCJtxRcPthAObTIn1rf6itY1zpu7Ot2G+6mg1fA0SsvYbxNMc/n+mIjScYgP/dau4gsHx
vhl6kn+IF6m3eG3T2HeOfD6bMlITgcgMrwRLRm8ODi2LfNhWsQUp/zAHwx3i6EumUrkR0I4pBGQ/
YH+tLATqhze/pmlCr/7t2LzibskoniVGvRfPYgiG8TigMi3ckG2Oqkk3c2nG4OnfYXCkjP3iniIm
23CVz3qCqaoGyaoVuLRE+SisZbO4QgCl1D6l0WI7n6CTt/1Z+hZfdO2XqG+zRtszX3te9xa6jvv+
TfsFma8o5y1OfSmu2geEpVQm0Qqu/hUnv8RowokR4LAFfaL8NjfDRGbgUTRtSoXYs9V0lf9TAig8
c8yowZDcvGfhu3i4CBb0oPElgRMQ4grG3ljwymHiAEPSkoP29NT14WWyJjbylhttR2xL7GPStPLS
spRcKinZl+UJUdC0RN2cGwWDb1sECLyX6J+tvFgif64XIWCtSh8qlvHAH8Pi1NQxI/Vwsgs01Z4A
M5EVJaKRgxoKNY8UrtWHN1PSF1WLe43THVUqDNUrNzKkAEqA5FEGmj2YEt57M3X5bKERdyEZfyd5
X5enUxycm3VRr6/jzA8706mb+b1Rlh7RaQ1/jYn5UcqX7mV7BCYTfLU72k81cKYKGnLIQUhirg5r
FUsksZZTUNL9phXH1uLrMiToW4eG+/vdNCWoRY6AJARgckL2unoMggh30JpTsv1AW9yGHk02BbOs
mVPhoGnjkfLmobnhVol6kT7mTEtj8CQO9X9BV93sirB79sOk0wrfXZGMimxAYD1nWyRjrS/shz1p
bjHClfhDiFskLpsBLU7rmAdorS+KsMIFWYEx3jbbYohSNGsNA1/R0yTzhChYlczrrRwpdnQ0gQEH
VM7pWyo7spiG6w0o6Si+m1KFDMTx61udfJW0BbtNCENJSZJSOa6n0o5JeR0uhjMHaWO4JSkKu2XI
LNYeYT7XxAcShznKJuvTervl+jSLYj1unw2s2NCn8HO5qIuCrEAg3LpedrahVoyEtDkEVBQD3kKi
glbVkUYYS6vKTp+ZhEXE3W6LLPc1oaNBNo6nEVI1ezbfTDC+5TALuCNNUtOjPvSNxKAbtcr3ih0n
39E5hjWV5mSNBtyygjRhADHccZNjoO16JEQXpz1/h8V30FA2mXAA34b0w+qdwyU1Jhd0ZaIFCQo7
u32yP48j19deodbGQxX1Z78qpak0kPN9utiTsBkrDqN9vtbIkVVZS/PGC7ijkYFIoAjPlZv5+Kq4
MbKPCDxkeL/Jx+zlQ/eJENwaIhTcxYiCh5Qnd96MIi4VnrbIzzZHlhzZwD494VjS4l7T38cRr4H+
m1seOASrujyA8uESloB+5KgvmJWYo0VdasP3Ocq+fhGHQrYAYQSwO6cBgoRTHRnxX4x0YT5DT/K9
GeMu+XlGSLlbaDUMrB7lL+/uH/qNSR86t8B47VMY3jZnr+oOMP0wCieiVGtHqG6lwD0mvg6pfBr1
1iPVv1KzVbRLKKBTGoPXNEVqnrks2XZkbuDSWo2ExHlCY47tX+eQTKgLG/L+fqP/ouyGLHp1znsG
0qSi6Y5Uwf4AGardtea4ETJsVk94QECDKSxt2wsaI0bMan0s6tvj259ZQkfLlersR9YEAevqaVL5
QYNgsVMA9gEHtJ+tQuWYsKc6FC3W5fOAnwHyPq0BB2X/rxZ5y+u49+PHbVwCvP++zk+9NFVk5dqX
FKhbwy6YT4eoy8NJuLt9ipJXPfXaHIdzAJy91fxSu49KXWFJEE2FTEMVCrsNu0m9J6sIpzzfK0s8
e3m3VGe3Ln5qyg4Ex+OzaetHKh5FNNBSrUxMgDoZa+lKB5R83rGllwMF13k08nErDOS+EGXZtJBQ
F2RC4f697buCKbCyB99xuJF8rnhYkoUsa0b4iumztl+sPoLLypwYNrpQpjX0xYARA0XAaXzToqDq
jQCyNdlZhe4x2b69aurfJYtd6m5w6AbAN8E4gPJNpviZhViJfsbFRZooVOl4Fs9lAZyKlxTeSARt
C0YQjvp/MsB507YDqOvHoj3QFxqS2bjwrsPowf9URUKsh0eef4AqsyRh/T0ZXUHF83xxMFIR7BP1
5iWImStLxlRMAWvs+gETC5yoltRIPz811Oyay3I2pQxFcKxmTaWctbT9c2vQJ1s3tFfvRVmgZUsn
O4qNbGKkp16vkRx8YPXNWQSv/jBc3/fvI3V2WopLeIb30/RdKv2efdvX9xxO4PgPBEayUrvHZ8vk
63kIFkdD+oU57xGr2SYKPt2bXbtTzdp8ABgdnkLejVv1jlFwtmrib8yyU1zA6vjdPGrcNyoft6Yy
zQDSmkVbGQjwzrvMgktZNH9Y5nm4T3hOcePSSiF8NR1N4KJ9c5kdxim7Riyu0enZvxVlskX8jfgK
6UJjblKsyT7vqD35yGvvDA6/YolP242QJNkqxtSGY+7/Lbqi89JesX5A0r1QhugKN/TcmC9jq8+I
1+093t54ABfYWjGOWqF/lyq6URHOMF9KLLRnc+rQY14m9TqNEsPQ3fQ0Arcu3wTwsrbvLFp753ah
6xwX+FooTe8PHrNFoQvdlXhvZwNrWg373c0//0LJmkiBJdXNM3J/tOnEQbE54s80zxIK/IL9xhKE
7WnYQWnwgypwmbGmsajWIH83Oc0BiFh1QQTvy77Q1d0wWhprpdZK2fKC86BtAluKOaG+zFjn+Wd3
lA92bX5239shODfHAifIo0kpuOAZZSCHbp3Cc7CVHUJxqMGrMl3dVZtGX3m69BhRWskfToMIyiUJ
it6kurzsUuE8oYLOz5LihCv060gwUIhWMoNngTLFmzZyC8RGb9BddXi/AtGLaPjKEr16xCBV0y60
UaBrWdX/0K/A80hH2zzjkDl+GvPCi4yhR+tAu0sVclAl8lK1EHsLO7d3zA4v4rr5Jfp7Sc2TOslF
IYhztTIQbKBopgvFcmtB0kTykwFrNLaCk7U0drF6+hGVk051CGgEPpihqtoTn52Fafoqk0Bf239a
HwvCEYo1Oh4L6kydy8y4ZSeck3wEPzviWdutKXy2ey0CiWyIRq8Uv2e/n5aKkQrp3MSwZ6JE8tVo
neMe0QR0DmJMxAa7ynhSU3tZMFCL8ap5NmGnkeP650rmaLB394UkwwMIBoMfymM/VRBEqiJUQeGU
Ieoij2sPWQyIpxTyxH/tczEevOhn42WO/+vMk/zxO0x9dcRyqLpvy6vsnsED0k9F4AXW1Y9P0OVl
J3cc2ZfWGNuaEAfZ9FV+k5QIULUwfYHByrYLlrDcu6WhiC7+y+hhOrMwA8AI8YF1lxg93xo8YYgR
yBtC35cALUD/4ylip2+V1PB2eWrkAaYbatw0fNqIupZTlXyZ5e65bWkug/7yvDw/xofhqJPloeiT
kWIvkSPn2F03ltKakNmoia3A2LzDHgNIplT7emRprp1wboRya+z2Xv/JsNacpgRYHl7GweraN+Vg
4NJ8SYrgfxECOPMvjR0Slckt4lK8SEOhyfA7WuArONCi7ikSKG8EotIx1rVj3bLlY2wYwhc61UkP
DLBPIE5P9BTrMRbpRUZrWGWMSzwM+JRdVxbbj/MnTdPVn0SDBPxJ5LHtjWnfWvqPNYrZ+PJmxmzg
HonjTB2a5WItqlKLIMYYIE5HBJvJAE5zsF2Ko6fJ/D+2qqiJSycGtjJXYKk8gRCq7W6NKScjXG29
/raY3vOFpPuJH9iuhIWhVwwYTYBElBMpwL2W+hes4R/XfYViSRjeRAUbzxJJb3W3DewdR6y4nw8y
0G/LXZh3nsk0DwTrAT7CtFk7SPgI0uMSpI9Zw1jIMn9Y/vFxXp2AWbTZ4Y1VuA0SJyUDE1SThd+9
NZYZVagV5BzhqgaeXtsZFXi18wRL2Qf68pZkfLIwFCs4dcSMnP9oMrXxJ5kNMU2qSAjmVUWf2hkq
Ykjxt8+mgyw/i3mGkpYmyXpI+V/h/VelqinkSyywO5lrZlyYDEl12kiImjzNN6aUew+C20A2N6SF
kFM1Sr4hvrUOrw2PjCxi1bDe/H1v0JWqiDlWjV/sXYkiUVsFaGzzEc1H3uQSWged86GtXFk7X+vq
BJhbZ0GfHtKB8bnu4UqueVFHgGtjeJiO0PsfCGH+EtYHLHclDQyTh9Or9j+GHPPFrbcozj5IjChK
FQzlNNRi/tVeUC09oktZYWmy3wvOw+NB7ESN8Cbx3RWleTenrk+nEdX3ST2PVzQxHhYQbIpsLyOU
lY9NpwStdCki0CJpEfdvQ1OtIGcfRO+sgSiQ1qpx0KaQoj8aMSQ43WgaxQU3+3mOEnWXhfqkpLF+
k6mgN9HgLk5Di9EjzIvUya9QSgKtzR3A7j6APtgWaRr5CY7mxQzKopJ8zL85oy9/c3jJnYPCIyYj
GP4s1LZoGm8jheulcI4AD6km/QLO60Wicbc7yeiV3Roy+7BB0duV8IFEM1onaYdwFdoNdQyugeUi
0Q/sRJjNYKhDun7N7NeIKyBpg7gZ30WEwsqHpdKZ9IlZwU2GqmqZUDDfClfHbE4wdWkxza/4RP1l
ebs7g8QlfmHJPHRuFLdiaGNDn/nUdJ9pjlRcMI84VTbiA5ATiIwrTJZKDKLUj76fDVTTkCVrUZQe
BCuVh08povl4gYNP/10bhtlWCsNwNzJh/W3LgFLLXK+apyqnOU4XmsJSKg/DQPipjGwZ++oeBXzr
qGYXajO67q7q+6zM0KnVSV2DSgkR0H+RN+NlIDNa6ZTNhZ0zUWfAU5W5jhLGlqC8XDkO03IAgFk5
YbcvZT9DV5E95mzF4x+y/BJHfWfs9bFUByW/nh+8lG+wcbJ/w8LS7+Y+jN1RvDwQ5G2Cd4Jsbjq8
sJK0RW33VoRq4NtFkeuVLdiG+nzQmYeZieaFKhCfvLlWRrsHcgHSEkzkrWdfzEgZLlOgEu3UqDpj
jybn0rdxHYpUghGLrKBrbC3zUGYEEGofMD3V2P0i7e1fzMY6+4kdXB2KDKoz8LGtGXmE07blLH06
nm0a0ynpHl2EbZBqKtfS1hDVyYhrToisJmsVoUG8rtr8pFAVfzu8baWA3wJoDVZXY3Ao9140xyum
s6aW5XHzqF+RB/IZ6vxNoHbbXZ37u9aQrwnslIaLs0B53vP1/O7jyhj05qkljhY4YvK+VsJCu8fC
fmQtFtN1U+toGHE1vl37ACIsCchsrH+NRTrn+/ioVznCJDFl9R8IeE5GnHy1EepcMDYAsQZyTBi4
m2V414YrtaG5W1EfxyJoaXMzmJzvDHSiYmUTLBZALP4JX0QG5sJjin1T5ybclsYWqCToQUtkdMW/
mnyPrmBmeyitZvJkut9YJAKFPSgM8UUb7fnmuyiPReKw7lvrRC0xd9dXGJBjkP5DxZHZ32HKb09Q
XghOpp9dENRXUTFxrSH45GxZhonJS1l3I9bnxdPu4kGoKwJjjp+0LVdgObJRaxTCsBHUqsn/Bz0q
PfYplx6i745tQ2q3u9RJOSFEeg/Qc8pRMS+6xMjP0F5jHkor1LNkxsn2FlsNkX0+49AmOTWdw9B9
Ar4t8Tk6/1K9x0Y5Uxw1ygkLQKHAKJEtP1C6AA4qEq7bXBVd149qutTcCMuVk7v1nm7BPNxQK293
j/sVlqr5JEAW+k0uSNQBx8U1taYogfSPqWNXaAfGS8XfOuvmonfSYCd3+HpnI6sosfTRK/GJh0s+
N1tRMuUsHa2vGoopYZ0A6TVymEt4mRO3bWw36G6bEYvtmWEEUtdKutD/1MGSANxvszyFFbXouJIP
KrD76z8NhJHG24gpxlckpL/etDGDrsJkVQlJZzP6ObuYmrYqBzRockmD9+q7krI9y1fW+Xh8pkF/
30rtWElAdAtoG1pYfxdS1eqaAhT8efSBHDJu9vVw99AFNXar+D3V5cCxr6fad0sFYewR0Pq1vkWG
+9uwg1YeiRf4RtMC8zQybj80x6WbFatiYFXoXlPhiWU8gyG3jAcIqxuOGAKl8/1DqAU1k4LB2Bd7
8B1fkF89XO29Cv26MRzF65o6sWw4fczw8tjLbe6vHohwRqSdLHrgJtXjg9QZtQOXDquLLsouvob8
55Ko9JPoA9Gl8kM5Ra2ehpXovNSOQ5FrYDHDjVOsS4x6MX7QSUVxlySHqGHMBc3T0x3GVWj2v94Q
CTDaNAsGgzkhHNbzoeC5pA8/2ADMl3fQM54w2Kp/x83iryPgBGtmSj0gON3vMtNb/srJt64ts7vy
/otgfGQNdW7vSJ+F0a1NM+Wo/H54QvjxFHc3TtrFsz3vd7ODeYkCVZ+ufaQQd/wqPnu49iCRSgJv
q2X8NYmnhTwAMfeaudoZaM7lU0NYkKS+d6cmigCD99g+Hvmqhv97hiKC9JbTPpG8kQ+HPFL6CtpN
zpmtAKW8JGoNYCjCL51PvIGY8voLtmkveSULtjRPYhyzN2Ej2VdADjakgnRCwDY72GtobS/IHW6y
6jH8E448iGzt9gCwYWTLMWhahryjOeWWVqrtVVb8oJ0csy0uu403zMNE6ZDHcySTsllmFuvR/zCY
M4UBbkP5+GQ/M+LJ/Pg2FaH9UXD23e1+pKuP36mX7gKXjk6KQSrXPnqIzre0to7dN2aPHDMAsgcx
8HkSu7GuSZZ9r5NJQsuFH1fhaPvzrGvHavZNMMd3xzRomVhl0kWaUXBPlcponxUEIfUif1mjbRBa
3jf7s9x5IILB2QtCn71JZNY0I7E1nMLeiEtnVjrU5XI1K1esr4raq/ex6c9pyxUrqSRtssY6wfPF
SjEPDhbUT4HsIXQVVcLm4sYMEr/qG0xCiaU708XoQoi3Gg0rYj6CsHMQpyzrklh5Vvp28c5lua1V
w2OXuyaPDmWsQN8RwaYNAOsxRxtOsekFw//OXXTMfCsy5yymE0M4ou8Oo13GjA92K11Wc3Tl/QqJ
1WtNtXdWxodqQiszw3HpswizGy9wzvjo17vee+4ht4KcDmzy4AGhHf94rDdnPrP58ei6Fr39Levm
n9y+SskyYpURJcrT7HcRCBrTgm7URXIT+Dd5EeWgA5K6weHT00va75TxDf+N/zU8/F14G8Uehbln
8oDo7jnTVbpT6Bp6lGIL6XEU/2N7snlvbC4JICSwpBCkwenjLTnaO2jHDSnnRO+4vc0bMMf4eW8a
9z8B9svBX2DGNKPbLwPRVhwLqnkzbYZ003ThpIxlEtU3reW3blGngnh79oVsJC6UOTDOoxFibaog
fUvpv00MLKFJTPxL/iQXORfKtC/nocDpeYIHaYF0O2uiyU13LKQwbdE6nnxlpKHp7BkzxSDKvhfu
9O/6QZPXTPPlBvYQxfse5cyWkeHjt999eX5v61EtSil/oArCPqYy2355pwOV/HAx1g+hGJmGwF5m
IF1CsRRBqc1g8rGqQ1MzCdlrWkKG9wvGq7v6TYl2Afw7xpZb/vfmefFagEVH/f2yTY2Vt1ZNOPjx
NzG0nSo2/2s87/wK2NFUMLRjzT9m2JDNl4PjbDIrF0u/ZNW893Vgy62ib+PAZMD4HKcXr88bU1jI
ZfBQ+8hZ3RZ/RkJwoe5N0tHnB2FeDuHOgJHg9brJ3TGF+cb+1pzWTCaZMQInySJRYZxNqhjhnKil
+Beitntu8wKnt7Pc/M0/NBSiyxypYsxI7qegnhD/EGTN9SZuV8Z2/al6/LmBPUlEX6xvLKLmwrNU
u2KHaOFbGGyXS6DSZH4UiQrlZ31nBDgNa9UGDnV9vLpsmHlieXKgBnENHnJk5KwjIP98+vjZLpls
QTOSuImpfbORbZcXezSNb6uf7D/flBWGCrUj2mq2KIFlI8WUkZfD+JKMTtP75tCwL/YPs9Hb7Afo
iwxCuv3KOfwU0XoU/Ad+jFnaxeFweWSNe3aOtKhEMSbmIyYrSb7XcoahDmsAmL7b6qRKfI+EBYe9
G+B22/ahCJPpagf92eeuwvIhGNGuQ4i1bQKKn4z03cChH/R7VSFkbTDeTfhZUZWFqkGvfQ5nKd6n
qMNkqhNEKre79ZwA3ykB6zhsKa5ruPJnA01LaVEfvZ/ycgRCof3wGRt0nUkM5A93jX4APxGhV5tA
07ThytVunmblKfTYQmeS2biRtFMTiBQkjSuNpdlbc+XdpY4ljx5PPW+E5ll7dbPNrulJw9sSiHEx
XPhCwNm0G60uyXk4yLNr+hE1cvA5BI//+qWJGf5FeycGSmNOGGVWvo/nZ8dnV4KewUDsKc4VZiSf
RSQnfZ5wX75tw97uwkKqyJ46C1mDlrNRWX9RobgYx1A3ibJN7xBPVDg+iTeEvnxYAl3KNcUUpSp0
KK6uKMn4f18esMOHXDgL+kVleXOzjDQOgSfQp7nvJvmK+xblKeaqfN14L5vo+yL7C03NS1Y1oIxM
5QmhhJYcl2EjhddYL3HNOIx8sYiWPXj2FCibz8cb/giv6dpCsjxZVVlAq1yxOxjQ/CrCsfapBghj
6g+8tbOQcIA4ttJIfazppCH0q6b1siT5wgxBZw3sQ+3thIO5Gqj+v5fbzDAmNIBAF1RM2xsKchjz
nTfcEQqFW4Ymj4T7P+9KNOk/UROysct4yMouFYUF+kTuaVlEKXgV4skNZEOBY0JrGowkRkUg7sEg
yUv4RwSX9OKKKR2CU2JMsiOs8XF2Kyp/fpznGFIcAsHfBgUQ77PqgwKgo7mI82SmUqyUJWDwdXAD
k3bhevAvXTLnBdCs400q5OWc7KVnbmKKWJ5290uoHMNwDzlRZOw0F/U/UJSagTb+2OohnHrqxd3f
X/8vq586rmdyNlRIv4rmzZ8Y+HHZJCpMOt94yW6Nl8fpHHfEnrHZA+rKJobohzKIAJ7KB/oZmIKg
c408Zbz4MaKYq+ztpRCkX+onJrSgxN42zHDPUmzM/I3LMpJNHvzass080V+c15jKa1wu5/vXBHgs
bzdYTj3aYN6gBM64iZHhK9Ix2KTfX3HAHw+w7OIXkG/ioXpFr5ruNreAumUstfMG51QMP9m2evms
pYS5mKRiS4iY7DRuPG7O6ALfUhkBRVmTfAbPgM2i+plxHPHtBPNvNEU8F6zpi0WgHKPbi5z3h0R2
RBicHcX/n44PZX1A1zpSiN0XSv67cTYT54D4vJmpYESYMFIlhwe1WACpRHt6EVCFih/7geMWBxAH
QOqJUV5DpnhfrqQpYDf1S6miqV9MQGGr2Oas5lwvQT7Z8vNFaStpxpA51vAQgK1edbIinUvmRwyD
tolTyTK1rIZwnLauxYslqD84U9VLn9aG9qSBdxfLEur19eljDxTzGqQ7t9jYQ6/EttMg1cWYluJn
PaP/+2Y5PRvICULqSYGCFNPyoBzGPoi8Gm2U7cK1iiF6jKBiGdd7IrbLXKTWHT8LXTQ6kEdQh7x6
0rjcNPiZCYCdHdf73f8zAOE6pGoZ1yD/qk8QFdng8hTYsdcgjQ+dJvhPGQWz+DqXHZ8ABkwNtmCj
5coF0Nn/cC+tyxodwXTJMzgEaskcsXg+NMJp9JhyLK9h8G8yejm7/59vc4W/Tt1egnNncaspbbB3
JvQaDugkOrHCREJ+4oMsCqpNufXuQ7Enk3WdQnQWGiowDeTYNdcKzEmz+3xM15QTZiM52LCK7JzB
fKPZcGnMxUkerebeoDqhV9cEXR+rw33GLIVKr+ek2QXujZtYZpFei2LluieystpIEPu6x6nnpOR4
mW+5YrQ/k1bU8IZf60DhQqRr1fFGfR4n7pqw0KnFGa2V6XBDAae+yzPwwWgcukcKU4aWebD6Piq7
yYfAjboLv26/E/ohkIh0B7NA3dvGJghjVAegIKVzuT54/Xg95e2V+pDNXV3N3/CsE5W8rpG5H7z/
MGjr9TAMvWwVSrGv9cW8zOfOUYcprKIdEcPKmoxB4ftrzLl3dfPKO6lQe4cNeQ7WJa7I+aNbe/f+
nV6Lq8r2c4fl7cWljhf4fKX9Ho0CgF0LtRc/f7XkecoCOTaKK0/61pNqITjNnCtJF1lLu6WvftT5
KFJ4/tUAmn+yA3TV39W36I52oTr+zBjoF0Ab07dmIfOvWVhKbuARz3RlxyHowi1bnq6RPSfgXXcL
3mivxX3BhmWkrDkE7/VLOG/mUBe1s1oU2+dn1me2s8N9odvBiJHF1MrLOJt4YznvThiScepBXRsJ
MZAQ+jHcdMSKkVqhBpSq3K9Y4eME4IqECaKAl7j4+vGZCr8fMjzY/mKGiRo1jir768d7nmK0irKY
MCWdtBkSziOkfehU0Num/PcNUNgp5lhRPqjeRxoZG9gCHTJlOhMNlHFPAISng3tjd2/piK3hBsoz
xqZ6rQCav8IU9qjM1ag7GiGyYu+J6Y+Ju7dUdN82dSYGh21Rp43Oh9yHb0VyjIAi7gxbtu9Dn37s
fLkDTNWJ0lH3qH7M8RXzI6Qda3j2PxlLpW1xNT8zECqmqOWL6Y47KI6zd0PX4fUvE+p8rsRi5X+h
Do4uap/iPzjszYTTVVgyq1JZbmEMjOAeO0zen1JdP+rX6xXf8mCrUpfCZqhHePfMnPuy+6RJ9FVj
Yj4nqMa6HKnxg6NrmowWjoLgpM/xHHFr3U5z9boS8EzQ7POvbt7f1+dPSCFvaA0mONvZ8qXJHK0y
xpk4MjjPQ2atwn7J40rOVBYWo1rnSVldZo52V3queusmzJUwy5LarHjtx+ly1lA1G+0DBPcSxRVl
5SNd/+oiyPwir0s7Y1eFS+oeFWJZt7DtbGX/ZK++Dux0e00fmzCdRKgT1HmPsStaZeY/OJXP79AD
fjk6/Ctv/vnPCqdamT9WQJvssJhUi02HdZUYVwJzcqEb0Ns/WjbXvM/SaJOzPSGLBWEdxhFiq3Gn
mh7cBDXjRtPo/U5TBERN1N9xYeNR0bpTFI1VF3cI72/8kqeDyoCBu1RF+kupjyGf9o+pSDYCXTMi
O2xm0QNZpezcgBOjZCIKijlFRySXg3xbYztgxdF3Kcid2xx7imYwxqzbpx/TDFxgum6oXFDcFYyZ
JNgkTWbr+X9a1HYOyzJBTr/XZ6CzzJOa4jbNnfxBAf5A5A5RL7SMUwRg4fC9IZNBMDFBMDAcJs2i
THQjJBHjeQJdxAjKjs5V0WIPABceJu/3iVqhugNr99jA6uao+KxRRXtv2I3AYYR+9pXGYemOe4F0
vlLUp65qp8vPIEkYfA05UbN7XSpvx6L+NVq8oJeOnrr261nRvDKLYf8pYPlhHwsmd/PQJQoVcOMa
OC/16LOhZ6y0FKOozpjARewVu62yxxXSSutBTYOKZSgBPHYxnC1qO7rfcBTDd6/LFt17ekIGSnfo
l/+yDpXDsVa6Q96QGpCTZHTULyMcPUTFDalxoPbQpgHddJzFRLE8/tVJjqJ0tvERhuu27QxkEJYn
5cqCHliOzhseTeH3YQSVJKNdOJc4eSPDKkum+FNjSbLyb53ZjcGCmUWUxYw5thNWEeQo3SDGLrpm
O0RXJdAOnLy0G+peg7kpAfW/WxpBwgnO4d5oScl5GMs7YsEuKmqRLZjbhA1IVilpQTMc0olTKUQE
4uWlByl/SZScg88Jcuo+Cym4JGnYyG0eTNj5g7nehwUy6hA6b4QhVrLXl8Rw6khygYBRvUAtRmTh
JhyrfXSsiBsmpfh0tWQnv4TQyFSxsP6rxHLiW+o3pcDH72M+XMDLIwY8/dnZ2O7+lCu82r23qNkX
fICHbjwzC0Bt6TBJlbmk9KiDVSGr4uzxp76t3M6f8nZrdsMB0cs4lWFaj8938nl/WUc/lDzN37Nr
oFs9iGbw/nPbSYmUMoefue+qtsQWCVksdxRkbDoXWzH3fKDKDVy11AFY+kxE0sRmQ0pM0Ijn1mvH
7kC2JxmDDYE7cjiEi1/LKv7BAb9nwcl75N5sY07hK6ZwG2wC30QONs/HCvFVQIgfbL0Hw62lL4ET
40cDvg84pFHV1ZhbOKnP2gmCdKQYJ4PT+dPcYWho98a3yw6FF3FIxkE/5/UTojiv5jtuf4iSSLZ8
Jw+TywhD9ojvstfOcUsTFp2f88MCtl0FJs2MLBY4MgsJB2RjXna7AEq92dfyTdXNyJUga1zjfVhC
SM1jMpF/F7E+oj8eaYNbCf0KD1qfOy2lO9MlKW9QO5Xsuxrc/hJt9zJsQNkbw8ppQuForK0EDNmQ
yG9jn+czOSkqTqPAD702UQNRv3gIxDtsSTI8rN7sKMR1cGDLUdiSsEorzaz5DsKSCVs8iO5Aemd6
u+W4AwSWZZGYm8DIhaR51lLooRfH6o0wakun946MyLlgMWx9XfZo8g5kUc3k1sLJ31HjAdJ4FH2Q
SNqJPW0UQNvyXAlfp0aNVTJh1YFfMsGr/nf39PYWIpZP5u7jQlXzkImMAtit4vAB6uC1hW6rVUZZ
Yfr0FEqLyVUYHh8SN/kGYQfHO1P4Yvc+A+W6KEmMEqwcgMMX25hiz3M2S3y3G/vBe38t6H+PlZTK
Rq3+IuzkJQmVVdEseypYbDx+cUk59RZNs+0kbMV57biABnwIbE5IrWgkknk/ZpBjQNt8pToOMxDC
oqvaZ4Wc9pWfuuyKjDxyyJWeTDqPPPHNSjBHMsiBr7H3EsEAU3G6G+JE1kH8bNDC3xVbFgiIFTo/
YjUN7wCz3fI9q0x/W/jqok8uI4m2LpavhxPXUWB47VLETgZXFkMgW/Fm8R9RH/rLTSXO7OoVoJEV
NbDplSmWEes+fg+/4aktzsRmJgE6A8JP786GZgvWQI8F7Fbk2ulCKez9RpsqUTBx1FfVxsoOxZWG
r91/e99LUIAt3ZuSTiezTSUYEYqAOQ87DpDH7xoqSy/cwUnLi3S9J4opxxKbQ6I5MQvS65o/jjNu
ELpRyo0NC6eqaP5/NvkxEoCtpIgIrY8ZDlczjkeWRj7IfjdYeXRInOwcvLnYMrq/sMKAUh1ydGh0
+R+GhtBizx/nrKwckW+IQTDOGbtaV6r3db1k0cRM8hYkpcPwoJEJp1o18obPURy7Y4ENy0oH9kRC
Tou/3WcmvFZcHwXdZQJPSgVeV5PqqOhX80Xfi6DqmFHSJqkm42QyAnUR9kDKJEfnIiDcCh5C4yIE
Cx/lvivBw8mgfsaCL8722Z0dVLbSRjiNwfEq2VODU67iDkWa2JUKHoGJc4qIs7cYD3MWMtaN5Odr
LnA80jmCDEjccw4J7kTN1BpQai406NI02xVrx3qUHIkpLgXHcvVAfz4T1BU35Mrk15yfPn9jNksg
/NRORvbHdKEjW6w5t6dLMO3bGNgdzfqM6H3LUmrXwdzji1Bn32JIMkHysXrvcdRMze+0w5bVUO8j
Et0KIhXrpDO0YJFovUUYzNkyIkZqIFH6RcRz1VFK9Pkd5PJxUBhyKV/nPym5rkP08vFDLfZjL8Bu
a8orDVDHb8oFjgCUFWbg0m7WON1kwf5EdARHEyuLYrdTLiTXYi2KIpm3Qem8IXPPx8vKnFNpl510
i3GsXLyq/iVZauIxALEvszwutNO0r1MJY4mvJcBYgDX+s1Fv5n8+h4GiN3o0Uyefh4H5KRu9HFOz
r6ZBMxAQbQGjzOZuInjvlqoGs7pweJvI8YBiedtDDlVoWTU+jGiN1Zg2+qiNB70te9L+Q1+YJpfS
pShxHfJBZ/pcFulHD54AdZSQeogvDj2BMbd90HXVPWirUJ4ZC/8UCT+es7sHK5HTMFdL3lbA8Ijn
PYIX8EzoG5iDhXM3hwrNhW4QNo6OuzRYRMolYcJow532SeJj+mYgjumAVaDklRpnjo0h2MMEkEpA
5wrn4+9ZkBwERTr4ByNsxVmETGaS+2GduCyf2Ccwpmcmqw1KUXiCOcmVSERmJod1dJ8MA3fezpcc
BG740GaxzE12IBESz3MSoaDw3OUC1ACWMGd006054MMzRM0Q2UwOsk+6cYWh4HMRpYZaH3Kv6FJW
qvYoQ7nFNrPf/0VqdpsK60WcYaahn+MRya5b5KBnd6nqgr4YnF4NbAeFkWxXyJCC0KiKa9o1DxeB
L+sYzqk2HmyGodV7f0h3LdXJ9s3pD5TBwoaMSGxFQUNGWk7C7dBqCYmyLX3UBY3qmtplvWLudXSw
WbkGCLQxVcFloKBGJD0tz9NMyUmjTAoWk9fwhALYqP/P8knF0B9H3eOrnmcLVS3+9t29ib4aiGmj
jLodkb+4FnaxFNVLZddUqKDMiub94+34+DBpnHKI2QFX7PcaMmSXvcnvnWl1tZ3E0cz+vm+Y6YAZ
0+DxYdV8sc3+49tdeV9CgjID0/Fzz6AXZsYI6jxkpu0dNYpHazObywvo7g4eLGppwz5nxu9vXNa8
uCJkotEzJWfPUXHEDzCL8+Jdx7QaAHAawqeJYZQ5bKjNtq2BpJuUydV2roOFBsPgX9LKeDYjnVDR
KLGijxujJXAK8GG7q5P7JVMjvhNP1IKK0U9EF8ICsbGBEOSpocXuiUd8oxdrlNV9IrGGjgwq9W/t
5eeRemk/B2QRhb4KAmVVr23UrpWfPCb/HlHYrWWSacNw2dAy6aMNl34Xl2AOit2zY9nAKtWZtV3Z
mm9yvOQ6tj63ko9XhH/rSXdOSSVxjwsuvRsLtukYMoB90sIzq45mixA8U+aav6cDmTpJ7bFXVy5h
+jj/otkxABt00N6/q9BZYW6pFl180I0ojJ+mcQEG90xrr1TQy2TT8VIbC78xWT/pZxCMsGm008pR
yAlil8yX3lmFzQZWENXBfzTs26Yz2IFa8P+DEL1faLjPHwuIoNR5H/kau088pgDu05E1eab5r1fk
7U22+kDvToJLqkKx/URCA6ug0ShCivlCgdjdjtJbugaLwbhAzdkQfL19KynlFHAT53r0yT+sjToa
aJDERJ6Ns8IHbGz3Qun6f8Ojr7lYj17QjRHLlhpypymwTGrL4FJcMXE4mtGkS3pIqiig0EDEKGkE
dwUAp4o7uvAoi9k7D/qy9xjiYcnScEHfmPcCN/+oxEKaw/1mRNSzil3W/vl1lF6VlaCyp+PI/B/U
M6TcQC+JMf4+T17HFZdroG1X1he3YvCpbBx1R8fzu9ACjPdWLZQtkgCYoTACzE26C1ELR5bU0PQD
EqbBNyWFfAxisABKqVPDnkX0ICeJKc/VDzrAWufKb0n3XzCuHr5TCjRIBHuWstGfdgu0pNWN4Urp
9ufZ01XwWx2JD4L8zwVILLp+7W33G4vdOT8g2xnpXud7ux/8aJM3zQeQh2ebaR+hRagwuaYhkqtr
htg80TlIXFg4xqlp68VzDABnpyWAMBTdheEzstmmW6fYWq5feKBnChvNw2Bw1q2zoWPKDk/4s67u
keMAIYW13Ema+7gEU20a3zuhpTTJUd72uDGHTCKMpPEOc/gjvNkbnzhYGGJ7QtXY3qXuPeHwL6WW
dF+55K/bNnQ97gIbnNqTD/2yxkfXhbrNdCa7VfeSFq/EtLk8+pXmPMtvHpqqKRt5hbVKOOJU+JAF
GKHfTZzIRd/0zQyGaFT34VqPaneiBtqYQgFrAG91nNRJTq+tuWQqf+zQu6/xhB7kbD5Z5ZBGZHaO
VKWJpvdizvoZkJ0rJsfVRWPi0vqgh7xzs9G6yliwAVJUGrB7OPuiOYScQIVGVAn8sPpZovnJeZdf
AephiIjEdwbyzN9eAvIj/9TBbkP/Mhmd3FC056Jt28fj+BzCPVF0QfGCxO077yTRQ6eqtJy2wMe0
C8g7nrkPdjJYRN5ZD89EYX+Q33lws5Rkhu3KzVxJDQFwOkijn+DU74CemK4xNTrZfzzrfqT4kJKM
TxZjdedhh3k+H1iKuIadptie8bNmzd+VpsCC5WfVSSMLGdILX2PKN7/ag4hMVoUuPMVFKAvdGK49
1SJYV/WTsCp2qqKhMgq80hUrs526USDALsTJI5o2yPUMr/XDAfp0Ioefc47K8dzBhWvOMn+eJXcn
m7VbemIM4FaP/iZvqHejlG3atHl/x6Z834RIvNfekF8fW58Xkgbqbcei3yyuxYKUVMSZpL7PWTPC
f6HH7/nzp1wca5Pg+J6kWVf/+yV0Bw6ptDg5XpCqKoGi9gbfQhqtbCnN7XxLnOYWu06kbRY3NRwT
cASSfwrlA2hr1d410SIt9/5Bj+UyMabvYP1FiRrRW/uahkgBvO8WpoRqYlkRNRk4rKJWoNiat6qN
y0YOVmvIIbkDJja0grc0ziIcfS8mXZlcc2s/+k4tQrFqdNTQkQ2oPg5Y63EiRpvr3HH4V4c0xXji
mGOmSQoroa/tB/VVh4iuAHbDU/7Et6vn7xZ26j/aZAxJdC0V/MNL/WsWLMm9Pct5Z405eUVI73b/
JTQok2+3JJPBdTWILla+dqYIllOnKmA/9qeacfrnlayvBLwxb1Pc2f308Si/i11esDboRHlkNgWr
s8xgc3cag8JMUFn8BxJLZ2HVAnLiu2H8QWyN1tSlN4MrUkiGdDtq1zpm9tTVpsltUtlpUX/EX58i
Ir1Tc7IS9YP9uXcwAh3jCmr+pwNkYteGed2BFV4wLf/0LmzzLYKaxCVpTnNKD1XW2E/Sk2cgZi01
IPBidIMax6kgFkeTU4Q0lrGVpc9qQIalZF2TSfq8U08uSKhKCytn8qMUdHrEFdyyHzSdtzwXAGrZ
4/kZ2gxyc611j9hdJ51IV2syM+DSSMM9fpTprTLIq9etxxIctz9SPmasPs69mYNttPKMXkmqJOsM
OAOOl4iK9PooeNHT/U9lk6vrkojtz6JImr+u6GgikN6cquXnLQdczYlzkI3iSm8kR9J8+AeGb328
2fu2fr6UBvKVNBpBTbJRw4BBDsCPqUWwsuTVfpxA8jX7ic1mEhm4ZlAijtj7EhUfDxh6PSlSI/6S
GdeBNwddcrrgndpWwI/STFtmRdVIckPi43w1wSK9dU4RNOtWUsXdBoYtXprneMiOu1zbxeQIUPlH
pCOhurSfC+TIliikulSudbDPIHCgaKetqXjtTt09ZB9IKC04D2TjPQSz+gxYCVJrmvdJcvVOvPPT
TI/+1PcK19P50z6/BIupde6WyYfykdf3xRk3TgseODLsV8I33/ChLmPx6bhVc6Neg7Cmw3hjBJ4W
YaL+2xMkPx+bA86irRH8fm3HmlJ/4itThIkvflgGBuskju+jabVHGcLWsRNEY5BEd3NX2va1sNVl
LZg/KcxnFA/4nmszCDu1ExXyXMJsH8pwnYv4t/IHhNuA3tyInDcllMy/0j75Pafo7y8HK9RYqRXr
EhmSRyt5UrhtCZMeR8qa65twGI9bVd5sO8NMljUqhVKUxVX5xQq0VzVnHYSIj0+tvcN9BpY3BxJE
BMvuiy10dVbB4iXktQiMlruGdH3rMWUdY9nEOICIuAo6/7l3Xlj2zRd4HclQnHOQlPdJuCIJ2r/s
viNg9lDSdagrERIJLytfysyuVxb02Pp535x4DBsFzBa8+y94bjg3SyYY+0O3rT2/FMFdaRCTVzTr
PtHGMHCKkYmS4faO3DybPDY6XWd/ZjYwCP+D98MF/Licx5KaZDfG9Gt3F5l2ew0QX1QwsZIkg7zd
5VEZDImaS7h1zQokOTqVZLLy6S/5OPlhhMGq47bpcVT/6s9T81+fP2qCr8r0szGgghIWzF2TVc0+
TofNVn5GrWTrqF7/nCLRjvC5xNlkpm3ax15xdcLHGfW9ts6cjZ8RgHmxOX4tQH8ys5p5vW8avpKH
wqbLPMeIEzUtrlK7klytniNpvX8cUregjMEk7NnrydAibcwJBBHNVlIUjXHQqncHpWZdrHehFHKF
K1vshlQIJ+dO4yIOlxh7V3LLj3dfygdbtCudmTuPFNHhkE4SjD9nNZxBPol/vr6wM3Ev1PyveFyx
Dof+2wvD5tfqDnZzLxGJ1Ct7YcKXAqhD9Mjtu8Z0cWUHOS79vkfODZuVqPmIxFN4ZQrwqX5URA4x
aqPM5QP+zvRitzmX8llH5n3L2eAXv+4ng3GIjBMq/rAz4bZkora7vdGIzOyOuR7gviVOSPcupNRK
RYB2nvztgLqlbaBrXyYIy0PqeUJoNrS+8ENiFQMPRFY2LxKHlwOB4XaEIrr7b2wJRMNXj+h5stnQ
qKvvi8CiOVzJNpIiCvkMeeDjMjK2d23J+Rmx6HWclsknDL95b0eRZ2Y0WkFSdqfXqML37kOY81ec
VSM8eaU65+g847mHip0h9WchcZQytEx3Y32YTc3Iu8cys2bK52PLlCl8MmVsQLxDVunlj+gH5kPq
Paa9JpVQlwLM92aeNREBRTPt4Ha4aR806FYvd/TLy9xywBkwmPKdvhipm1yDMQqz+yqQTVnZNeGO
hzC0hhiprzD3YttbMegVngMaaLoFLn+JcrDkftJKrertUWgnNUeHfaTzOfQiuliFaVPoXhArrLE4
G3pVb/eYPWrDSQKbDFwuFK0dwovT+GGqiG9S0ApdOXhoOid6bd+lZHV545ZsKT65+PVaJagT/u/k
mV28QbbuHjuJ6zOWsXjDrX66WN4v/4fLQw6qatxXAsxhGPh776aHzPo80VQcmimjncvl29NPSMOY
u0voqwGhpqHfQWkJpQuh1X5UOqfv2oDDeDFjjL4vk6PrzbyiT2Xqf22M5VvYcJmtsP3iWAbLmhup
mEvBhCkA7T28M2YZLKP2dCYSe5Ky71bcmQD8I19tGG0EcWXGy39GCyHNyqddXE7F8DzKAbmDTgmG
REPlS7eFF+1v3tt94vgLQ2v/bSqPf8xmFJojxz6HN66zTGRC3PGpjz0s4VDwcT2mNHwPF17AyHVn
Wn9t/8FWK54LdINPZ4MQmdbYash2lf2ePZAln3JS1FM6QE7qBhR4W0jruTz8UNgKUzuHGf6tKOPJ
zEOi+BcqRsnFGiKyuXBZvX5HrA+8hVFm07VeZOFlMcgsj7M2uljkgKnje/GQk/pcOdyB2NjJ7Cww
HpuXcBAfCxKCFnjyGQBoyqc0QUMz+0OzjARiKVbhwpjYSmWNLRSpV+Eg2tuETqSEJWN1BsnkDnwD
+YGmeVwcgI9RDCMWvNrLYIdeKyUCX9UM1pJ3IVc7bgCIZ4ckUAdAabtoiL/hY4t1FIBDBkHLOeFe
TXtkH4B1rIvCvHgoPRcbTblPGWClQ5Jxd9Fd3nOXetCf0Fp8JelwPFk+5xbeYr9mE5StIu760ytv
5GVWRqWH3WqafK1KqrNAvZTTdb7KlBgtYp/NrogbI1lhDKFi2rJ0ouAAbNdsLASEKqxIlv8kYzj9
37uZEfyIbOU2H+vAR5dqf5tKQxsryNF5E0Wo+JShqgVdDYY8vdjsWx89RRBba1C8+g8p8OZHw+7n
WTPC/JY9KVTNsvFWBq7ViNWISdeGZqdipcXWAYi+mkzcLmPi1XaMMVLqlhZecOD3HpmxWTpA86Bq
UJxN6RhG71AOCur22CMBSbugPyuVEItEA9YJUMpeZuERheZAs3zqon41bRvs2yXtn97uB4uVGeLT
PPqkaZaGTu9ZmzB0jZBQPV7vW9wF5tK21c+xat/NoQshkl/l5TNufo8kgq22OwkOGKvXmhT1N2Ma
hNz6b8wzzVsIZ/HFV46ncHqzAus0t9FrdMoxSVGR8lTbuyUcm8Kqe0vJORzAa78N1vgVYL49+lva
RV70NQVWgzhzFx+YmQKH8Fx2YMuvzhpdj3wgXOmuKVEeSC8IkV/wZjs9NDLI524OavGRsQIx74ls
cAFgFy7t/8OM6fNzd1Rn5O+RzSQ2+Zy845t051xh+KlIOsEMouircB8bBjf9eoUpU7Co4RlMuPBh
9debhLYidKuNJ00GRMIui2+xu1KosZ5BJjC/JmlWyJuUCXhJNTx9MtkgUItb0GzP/JgolYdPjbKb
11z99w0tmTb6ORrJeyraBBUoZ1pUF2++xxFmNnNYamgpv63XvYJndDxLo7Ej4oUToKkKR5JHyx4i
9Y2055Vtq2bN0tpLCMqWXZ2vaRg7DUHPvKidNKHGsCo1WCbZqEVNWWINOu/eFBvRYetUmay36+wa
21ycE82VV7oA9RfuAP396G0XmgR1Nip4bnHIhAMM1+8ASz6SzvClLpmnjVjMHTfqFmsdAbqd2OJX
cWH6wRBluIJJGSXeNDZ1VNBtiBrkokDZhMzGLwFH7bBDQG2tX8A32Zc3Oi2a2b/IGp71+2npGW7e
/bj147BC7w00MgAmNygrRRBkmw1Jqb646TsBJb2bOZzqCIIYW9Kmxf1p7AjtJDRatQTvU+Lnd+Fc
ni+EMP0NQwju4s+FTgoxjRp35PkrUrwpFLC0wJyUMh5VoSJBpnKYG+kvqGuvki0/CcqjhwJ6d2t2
9EfFo+lFKkbup5AwyoyvpMebTjNAwA1JfnwCJsZ16AEzd2XH7xcSpUxY4sRNcfGO6QLxGb2PkRbC
gSxUo+KsCkXrE+t+Q38vShJvk0xJV5mjk8xmDvGMfapE5OtnySLfuEWZkCY80S4GOTdgvON1acqq
MofslkNft38Dvw/SyAYLH+wJ2jY6wGTl5h1eYbeDEF8xW7rAcgD1em6G4zk9qRJ/Njg9/YdzUfPD
hGPl3+1NyTvm2CD40UnttKPLByoivnB4Q+A++CyQJ9xg/da7zTPZ98FCY3JO+0dnyjaXg9+3jIGc
g/BjFubHRNCf0Ax1VGexNywhJL//lwIKrJVF8TSdwosxEy6KZSqNkduEJEkwkHVyqH8/YrKwAp5Y
tNJUYSBtHAe0u5/rv00rIjA6oEnM5lpssCh4zHyRJHoswGgOutM3pjUWgb2+qvL/hqABPl6CbbyJ
3KFD37dY/yUQLtkBxVmSVtH6AsFY6BvbAiC+2N5ejTBxwOIBTOvjppQS1jzZfKdO5j7NU03kroQH
IkrzAjADUykSNRlsl4eobi8h5i67QlVhNlc3gZsQO0lExRILXi78W/BhHUhPZzkeRkn8uQFAktlR
UJ4D1++MN7eXBpixW8Z68HE+4JF7x+RF86aaQHuQ1gExqNxA6RjitF7BO9FTZ4E6HWdVmRV+uad0
HzfdZWzKJVWque4mxBZv26Sw7aMVtJRiSSggFjPBsfk94Ky3DObFRYqXM65v+TRmRLLUUD/t7JkY
xYONL0lFhkhRtHNHQJUSgB35kZNPRlG1pcX6f1csjdZObZ9ntkjJlaotvf2Q5vd4LzyRd/eNELx3
Xcp0YbyEJA9yMfhmeU2j4VHwWKFRJ9j7hK7dndRqn/fvNMKeDm6YxDhjXrhiF1d15LMX8zJAFFZO
KPiSYvw0BnbXf6FK8cKjei2QVHgRWFf8E+fHC0rK5ya11JBTFcFRWLwKaS94bWgWg0TAnxktmhf1
iBhfE35nGR0IryvNVbIbqF9KX5JoJG5IZXU0ZBhy65KWUo8gselxnGOq2/8bnmtV7p16VAypAjG/
lDF2XrBG19OY3LtVVhB9TVjvS6zkbDWQIl+dpsIQE/1O4kiAs0c0wjd05Rkh9PhUey7rnmSJNKyp
NOu3rDoIC6gjqobwOXHhkurN0JMVC+ZkMRvB/hw9w7yHTQa69M5f3q0uwX+N1rX52u4S+vDcDXfr
LknorAfOOpoyjcX9sf1++JwQfHhP0H2sZQrJwC2zC5e6wyH+BdCP132PC9AEuCxLzAjgTBs/nExb
7sPyExkXfqaKCd1Y/vlkWkpkfrARc06lwjyr46Yue2lvtVyTH8sXenY6iXKTmv24S87VVRBCdXR+
hbeEea/ld4T/mo1WC7mCWdeWTojTvtq2E6v2YMDzCvIXYRChF+gN9szOTVCWpsxwqAg/EqjU1jUX
q58UP722YWCezxJXlHEBX3PNLyluAChScNL/a7lodZo3HRAd0CC3QQju3afszazTMjYJdO/X4asz
1rLDCfksueUBiRIp4G74FrqHc+RZNb15aiYvoA9UgqwjEcYtrV6amrkio2Mzt+75qEEpyx41JPXx
SCO4hiYplVH5SVJHGSWVjuWcdCZf9HorpQpJ+Bek4DTwjSkvWodaMaP97XREe9acnd7ql/dMKk7X
6jBDYW60HsjxTphd9JUI8u7nxHgY8WRabRn6ldVWUOZ9oLuckVYeITYY/9z4s/lMt+vd0at5MsQV
YH74toPdw5Er0alQADY4kLEMkgq3+k7mHTpopyGxxiX9PM7lt6PPeg54yVDJdcs0w7LCEWe/UoQ4
M9Ico2w+BomkHPeqsYXH1Zfh0NO22YevyN+O+9vn8utuZ8P4PyCEsFUdvQIwf7IFHIwyXzArbz9g
xxEiVulW9OGLQu8MOADl5EI2xWWuL+xdn75PEWM4Un2hL2YTuIuZzmFhx0mMUKEJ79ggS0baB/Jg
zjZC3gEt9OjoyZ6x/vSoDa6TMFgevqR3bRmdjWsGqqZAmB++vQqtGlxRkIhNO1GQXJOp3eNNYdwQ
XpT2vkLItHaGey35TIedl13Mazud1X2u8L63wN4amyacbIYG9HI95fDcbylKS+Qo0QgBCi/LbYry
NGCRIPDiYzhUk33shRIRZu69FhrZQRWY9pWk7IGdFVc4AmcKc+AoYzYYy77SkYhVmfscmExto6+N
P+Jqv8tiZKHRuIT2NQoir4eiZBdXryhQTt5OlWEamepIhub9wk0JoaX/a2fR4kMFBKEZ1oRwZoM3
hvK951nYLmtW8DVvsgjGhUdBK7JapQ7wSH9SgFzO2yfBeyENpJGqWNYczyQYQwoZGRbZiMkp0cxG
nmg+oy2YDjuacF7FdZl3oUzNIY3x3mLH9J70H3sr9ClCAhMifB4D3dRuds8y3t+b1+jVZhsg/Pia
lHv13oLKHCqmTQsfYzxeYksE+QsJ8oMFRBfMkg3f/6h5t8rUHh7KXwjqf3VmC6XKl6ySVuDeOVPq
G+xkiR6fM18X/DyCxgcrgV1xtRYWFLuBaMrTXUGbfez9w0bjJ9F35bfwG6h4t0pj0cORbsT5Dc6+
L2fcWTZQp+hvGaED6snHov/YpUjLmW77gBXb+qHj+ew/tGvsD82jIW8iJaadKKMpvH4Mvp0t2Oq/
GR9IENHpyKqWMsPKgOlzyIGcr4Wfwx2CcKjVmdCbvgYRgQaoBF2w77SA5R9l0IvI9s/kTEBTUjCq
vPVXsRkau22JwoJQq9cwIjuBBxw/H9n+2WDoVDffakbnwCnn8i1EyTtWZZ9N00Y9s9oOl1UKaH+n
owghQauWU1MQvtkgBeIb6XITn1Wv3IYEQx0g24Pm51BTBc/T4v5y1hQ1hxNU2qalaJdHJ+yL36O/
9Sex0B3CP/lw+ZI2FXxi+Bg+RrlmDb4JH0i7HF+odX9tT7ywiipALOU5KWmJCZ8oKTeJXom/aHiz
yUY1/Mt6q0YTmq6VUiQ0aN8gWgeiekjkp2odV8XWSyUEeackt64v/xLjI5bwfrtqcDXRnxMNVa9A
W6ceDuDac+P0xExJPU49NhUYu9iQeoWwmsi/Lg6eYwgPPgPxHtjxL7sDznRcFvRkH1hiRQ1lAxvI
lvlHhUQHmcyVb+r42UNHDjLBxVBSaHP5ADxK/rz08aKjenaj7i7FVXUPwd7wrc1e+mpLV409qrjm
yOin13QjnL81ROoOZDmpncTcTgnRnrp1+DC7Vcx5S7RB7kdKkG+rfKRSfFpQ0B947vBn4NG+vqDK
zEFz9TCCL5l3wDjpD+iopjI8oJgUOkIuJVhtWDwSrtMLpBgc4PYx4y0lKSGu2Zuh6xGRzIMrmINO
X73ECqEY72WxeBqq/YzyFKP4R6+GQTjvTcn4+1tbKa6Rt9JJ7jOcKUdchpcCW4RBgUNOT2sXilCd
qmnPYFPuAJ48ZqDsGT69VeEL1H8OvadZDzhvMLPI+cAQ5DLiyKgUkrs4lYoJptsq4mp/+mfijH50
sgyjOGjYn1IYpBnPzLXraekkdinRcMOG7bF5HTiTmVhd7KFhc9P02LYFMn+F2S4N0i6mgRgbj8PT
Wg/78DNapTrwj7ygXBQua6X8U7e2i93zY13ADHRvb5oYMWKAO5c+PZnpVbA0PxwR8u2GswgX5fA0
z9q/IjofmNQfUqM8DIyz5JRocm1UkS2qhaKgW2/75CbNA2VHdS7fq9plSTMFh8Z+DA/THNRorQdO
TP+6ZizNTIRGmyDVSGiR/c4D6cazsI1sm6VXpnMVLs72pCikU/Xn3gkUkyOy9xS0SCqVo+Kim+qk
/EezhigGRz80phMCsGp/ZErt5IglfJ1vV5kb3k8idQku7Jv86vcTYPRcsGoq92LhZVF20tgW9ypN
CqKQdGjDUi0qNl2/eRZ8uKquRA2VpLqHU98N6TZvJuu9e5GYzM8vhKH5MofsEBWmW3hctULaJNDy
0j/rxgm0m1nS4D4fvoHWCw74tZk9tBCY6XwmMrY9Hd3xVk8cjrPDQOGG9eUOfI+1D5/tPzxcEaB6
Jrde6PRvP4+SZcPrXqV+iV/0KYfi/qAKgT1o8QoDH0hwY0EYcY16JCAPQ2EbDF5J94wiB/eTsJSp
a3Vka+Ws80oj/jW2Yy2lFA3+P0vGM2W6OldG16LChKWFwWVmn9esmnWh8oBHQndKQAvBlw6iCJhd
7fLVfZbDqB+2q70g5jyB210r6EuBy9EnM64MuA+lT9SyBLMuE7V+Ldk2+Me0VOJCkghv9KHVByVr
ijNR2mcwV/AHsy81U8A56eOobBmzU50cQudSPR0UiwnadwSxpprUW+KcU1dhOTaQs93irvUNekax
6Axf2IpiXtTXIPmmnsp4cLR6KB9FI4wK1J92o4rnSeWTNsTJYRN/1bXayB7ixvlhzktyPqoZtyaH
aycXW8LcsbA7cTIRikGHV+OM+0AzJzJFUDEvZh2bRPn1hLBVqO4AHiiIqYXOVj4fIx613XeL4AJx
jfT9hMNwde3nd5ClmLOZUc+rjwz7g8FaElbkjUoXTs0tdljGLjc+ERjFoCciOAuEtK2niIaO2dda
JVJYR8I1RaR9vbed/JZPi4XdEgqJ7CBfnZeCq5/HqbTOWLkrrdMInD2THU0a25NtshQ4TFM1fU61
xspLU2BZ8rOIMILneUy3h8AZ8UIUd+t8xjwWCpLJG/esiTu25SdSAG0N1oqcjmtUoVAkgq/dsYMi
Oy085hYyI3BMgVg7zRMCOSrFRkIDkkWQ8u0Sg7EnbQtwveC0Xk5Gf+FimEMDvkfz3656N4rnbIvL
JgROy3aPn8fPUk8eZPbjiG1/tAUWhwzFgEEC8OGb60gxudKtHM2h3OfaRvbLpVlRMJQeaYzuQ+cv
k9WGAKRXj7j+Zrp6f2gYLVe8qVr3Chc3pyi9pKd4RTyIt9E/jTO/3yaTMCitts2ACi2Z5S7vpKEk
lWsyv5T0G3yHCfg/7SBQxIbgck43SnJrgk5hs/qlMG8ja5xU8QrKq1BZOvc34JiU51OyVYDX5Vhn
Az4B69dPqI1pfkmsRob0sOdxiWs4GiATw33CnX0DqZVPHjWqtS9yv3kjCMGYAcjr5AoolUfolYRz
i5X72D4WrbglQa+BGZ6U4pcjoLv0/WpjUJgAX/2O2Fo800lua5RJlcW+fHAj26ufrNmgNeyfaYHc
pUdm758oj91EQOkzz2JmtXDPuy47T0sj4I1Ta2hsbOjTz6rLyy53eeu2fw9FCNvZZhI5dJvHbUok
MOV6tc+tUVRqBvlY8Z2IdConIueWXkYUX5qof9w5PgJ94+O1MyvGNbK5i4f9BvvUuK3aaLW64Rlb
jsDRahuAecT0MiQAnU21e4tU22MtMlshdwpYUoI+7VT9pduwqA1iakcFnm5k+Zd6vCDppi+5K0DE
tDstoKEF/Serglg1wY+L+ZY1bl7yVstXRYDtfqxLMKUB01bpR+EBWDcW37FzlMmMgSHhs8/Kcdsk
oIhmKB5/4R5nGh8S5qU3xEZ5VdOLNYJlcspNJLsjXjABWWyyl12G3I6vdGgWV73EID0yk3n8ITew
FJn1ak3ZTmQo/Mn3N+xLMkI2j3I6xd+AP5B2nZx6XhS7JgQ7cyvpjPKaFDGW2BnXlCm08KAMdM+3
nrfwygKntegZdzdMExpiK8L/cwsVa88zS2dASlVRI3t15AxfoJnDLalMJhHI00b+dWAFAFjCUSBg
l6/uX9GdAWgwQz2DR5vyx1hlC9e+jTePZLF/XEd7Mcc+K/doYrGLcuL66nFxmxG5fUtzBnrCTcc9
h/uMphP4i4q+cWFDuuDTP6bdKbT3qhdfBq+Rr86zmh5BeeLe3vWS9BSo+Ir7RVLFHuorMKIC6NUd
SEAHqODWXk5EghNrFonOnDSLfkLwX1zrE3d7JhkUxC/iwDpghmgVcNfZViAY1N9mV2TPM1waWIfH
x9o0cJsw/Lrb2FS7kZi23CIKQpEm18VoxzBbt9uYTQ5pgZDf0fuNNvSCtoLoLmhVLsXWc1EVfH5I
MkEpSW7mTMBSQKF563CoZmMzBWiV77CsnEpCdPj5H5uqu7TgQ29wBb2jOe1vuiE9HxS3ycBhEodx
hpPSfxfHfBdv9b3rtgwvkeS5r9hFrXS97RQ6TwbeZzyIBqYBiQLYGX2Clu8kkzyw1iUwD91djfgN
cEV//hXm1RxFRJfqpo+xeqvIqnxDW4bZfNYPVz5FQk1zyVlC8kXwWK5LeL2XG3QLkFcmNyJ9QHSF
N/jNW90/eVQQDbIy3aD2vxSYMCNJOMRoxWf+hh7swcbMeuhEUIzW9CtXkzUr18xsFPa8aV26KWBU
zt6GR+YATXuAhWvp0lCqhPdCyzyVvQeHbutgUoBLZgzoUeIx3BMtBklxq/hpZHXMU/EfwAKZK+GS
90RC7QtTYYN5Kk+JyHNyLYjNoKTydJON3DzwBJOLcQOZk9zVY52DtxtjTkiSXLMEbAjaua7qHYce
TwehYdYvnKsBE+/NhyQcySOuOQdTj1qmjdL9FGU6h3QzrVu/oMakPK2bO3Q/Rc3bFM5TNEwX/E/R
7VIGXuL1U3lyCk3FcQUDJUK01e9n0cPVdqGjmhCXyWdWPpx/axLIFxibKb9MDBCpEa7wHJJfxr1Q
X1cRek4Wi91NF+bWRQex4Kl0VeR6yGdtJqIajJ16FKpXCAj3CJTkovoVR9A2aZCQAoTr5+5o8wKV
6HU3j3HcjOEHhaQH8GqIvQnIDafyCd5Cp0Iun9FjarqRRPnxY7wj59e2OaNjGV5TmI7yRL6Y4ghy
Q3Egz1mZokZ4j0X3Pex6Sbw99UQLhg7HfCMadEAaMNT6ao3DALOUnUiHr9m3xL2/2OdJtAHBl0YB
ttH6BHmn7mzcTKToMOAOiBPUhT4PMRroS2AsS088spBG9SWW8IC4p9FheX8mIYZ7pXlP3UyJ3RV2
fBljX4GbsLSHI6Q8rFby8ym6BSGYIVueOWH1W83HuvhrJklTJPhqc4hlaPQK2eoL/g4EEr53E4RT
VkktnVPimRuIvMTXI65Gx5nIkrNj0ksB28bEZetmtWQ1pk5jVSS2ftdw3x75wmf2wCQPmhO4CvCs
EjinllTONnjF/TfYNUrn9WWIpOQXrY3BxAf8CQ3rXkTCdORDTm/PlBGCvyGHldIrEF3ScbEKJtRW
R7WZffQXRmmSsE8N6jtLNaHm0XfnUzMfr1ijpItxPuNONX+jilH59FTEfd7EtexuAjUiheJmhLNJ
9TkuraOfbxTghUS85nKucsbp2BZ7bnAAj6X88mwVXn2+97IlpfeVcG/LYgWOozxzvmjbdtO+3/0i
PIRq79ScJp9Zxl6zk16eycChDR10vMcDsCU+5fpk03R/FxCGnMI/ysmAtZC5YAkIvDfYEtDeeJn5
OB4fYSdhCHNi8ZfR8jEWzrjdsrifJ5OTBwpO2TuwtKMhamQps8XQ3mMOYwOtjAp8J/S9abFp+HEV
v+umw+cwOjRy/hRk5RBuhy9fc21vZ4wbf1J2W4cogPA1YSjSxbP+Tqv9CvDDf0aWteYIh7r5J/b7
oZHroTLOxLHKVI/aF6s+9fcL+nVjs4Sonammt65ZgjgKwav6wIBY8VZlt3VO1fS6w++n2hPEsjOb
8+S7amDQJrCRCwLcTnYDpVgJLUF//ZDfQCtGWveE3TlLdQ4b4Iz72NDTxEujCpRfH7yjHeUHbaWh
lmgSK0rRtOY3Xm/4xHkb9intiLtBqlVFoU7twCuKDhvdCl1WwWahHnKaG+IhOLcC981F2uUXQqtJ
YVo4aJbOT5dbiSqdygOoQebHwqcAdEgrVD6bDb3DK3/4nCZ/ZTKSJc0bkFzLyFvrGq36MBJqUIyr
CePPM2B5FXTQ5khkT5sPx6AlW+pV3XzPcR4Yxlc1p0oUKHX/wmup8TuXFYpna4aH8HtEM1lz7qT3
nsg2nY67Mu6KNtIs/Ov7o3nnE8W1fC1ZJ49R7OCCFFRi4FXxOQJa8ppqRF2oWjs/M6sFNJzF+x2D
cpfAkUZhTdmfi8t5dLeb9OdtSptYz9udlHPMiErxO5q3GU4k92lMGfA4QY4f6fGjMBFewwgA/unM
baqVCtyQHXm/hJD2g91WDFZyp/5J/NYlqw+XHq9cRJvwbmGuj29WJ+hui9Q7PSWOVKzxoPs0qj7r
hZyq9WCc2gjxAk1dY6uM6B1jEeJ7XcVw6uwvMnELYaiPEn8UHg6OoziO7OL2hRLtEx9ughxXoX5v
UJKF0Nf7PwVkgyO/6QDuxMkSpkX4mFufKaFbnRRjiVpGWVYHrDkJ5wDiBJz9L3kr1LFFJ55K8ffO
KNE4NxFknV9d9+fJceJD3mIdwUJBszY52y7f4fwDlghQ7g3utyOkNNoi/CHsf9uBZGYAxmdcTpF5
OMQmBb/zzueTZgWKVJzIpWfkMajCtzzyHx5Y+AQ+swqQkbSKLKSctOyMoNZooiPj3V3hv4ncWvzc
3cNPDJcXhKII2+8kbI1i8FX2AH49qQdNX+NVwKNcbPUZKkdXKsy29/uBSFAh6ox68idJBKEOcrOf
xM2y4CagNDEGWxRI33oLI5dNyd5Jv2Tf7BU+QYnNhIHHGKarTMqtJu9asrhWwOYca+LoQgXpiQ71
0abHvtg0SaSGVaaXERnlHr1g4rS6S0xZY5ejnu+BVyrq/2VzCOltJvG4dZEei/gwp6PQwXxeic+t
+0Iuaew2BcDv/9SVLnPO5hNB0iQdUtO+j/z/lZJNfHC+8wO7S3r1xLSrRgUxWIZRmOR5A4wXLhdz
0bsu1Rx7xbFpiGOfZ4p+qIWbVWv+m6fOpRbEtOIqo4jYRC3rDzBjcZFdLO6yR400JJRxmfgoiX4I
oGAFMZkvtqVbjHETf/dsdxey6Hc7f9lgNAA/eUV31A1daYHaF9JcNe42jT9g2ycKOwuPHFyRkM2o
FM6dcYfQqnOU5wtNcLYqsiBq1pCIcRheS5e379/ED9AcgQinsTwXZEd0kXmHYcFKasIxTtWdvhax
/PtKEJFjPw3STgEYvb7RbrMjJE5In0exGP1iJg5/p0dq7Y317/0NZJRpr0RqRHvDfLiLEIEh+wN1
0kLvQooRAqgPbq5Ors0PQW1e/CEbJ0aifeM6rcCdpJqrE9oDv0z2z8eFd8KmVwIcs1p9eTe8CWkT
/0n1IFm6gkYVk9SazeNunnPQX8wlIU9yW4dYKhcJvDLqFRW3+MlWgIqF/f3G2bEf0D3YHudvqU/L
ecyhQwKz7gTaicdYm1xdTiOEmHHRqV05OfGLNEnPe1ttf45W9oZpYY7xe1oD9gdOVqwxh42ymU32
Gw8m9zTIDYVcthaH5a6qDhCdTtIPRWSF3yNxZJg8747eR+LYzBB+xgMToImxphPu6RX5KLZJXQIu
jnut9Ff0xb8ClLEUtzYl8E6HJJKywyetrmjC/+C8LofdAoPzJAosRAaQgoaBc9jxwXV3Xl+Uf9q3
an0Dw2Af7abLQmR22NEXdykuwKm6ESPFZRYr2EDR6adYHPkqc85ziIawl9LxHwN17nx2iUR+BzLM
mnl6JXjMvezahI7pZLDnk5J89BS28DW4KvTMlAAhcTWefC+eh1JZnGnJ0yNVixY/xJQWiv5AxxWC
ZVx+HFdnzX4S+Av8ReD0fhOvanTajxx0hQfLHsphPaDlLghHYWr7/q1jhzVFLv+S8BuB/4kx3E8P
/qRYHnOnbBfHJ3jodjJXEFYxjVPfWcB4+QsH1juPIsrdXaPVG4mZcWgMbVPdNv5EI0XGTYoPZmdS
0xnCvNqRt/jKImwmxbmFBVfq3gxglmksGwRV+IfoApAghd+gATY5FzH3yTRLDSC6X8dygHIa7QiH
1Ggew7j8Kg+tf4Hr5y8APEdPrEB/ckhE3ihyG9KbhgUU7KAUiS+y+XGsguzTuwGMnbxQXYQP90mO
1lPyMQ5poGldxwfse4km0DC3a5VKaFkWR3z/e2lMALhJxiDQHeFcgVCpD7Jht+2nNViKM6LkQvEa
q5Wz0+ONv9zCiplQNu3bT9pFiC46JWykYUNFkn8dwgb9na93+XJpfvsToNUSGizgz6IzGmN8vgr2
l2mTuVkyDc8Ziyn+sXbK5lL8si2kYwUy9YyQ0xzrsFq+X5AQHRGJXenHYv4efNmbWatxxtKUjdqs
Enx0EPMmnr4sPKsmbKWL2oot08sIhZQH484fi9OvO77rOYyRPoTZdZ8VJcE57ZcZp6ydCQae8tU1
evV64u95E2oQCt96BSrJOGxkxFZqT8/WzTXueiPqK0XT3yWQCjlANCiyLi3OIRdt3KwgmuEK4vBV
M5pHK5b7lbnyNaNsHg+WCMXL15uM6dX/E3jfnU87yQplPbTnME1bIB9NNVnxiswGpogDWdXY0LK6
5E0Oh+xZBvcFp3VDVlH+sl632XRHrMCwFaeRHkuj5vOmetJk9I4wgrpSbusCQWl40xHJf2lrc7QG
HGbzCigCpRYGf2e+yATKo0VHnMaK13RhOL08rSp+q6fo8oee6uX0pOzd4gq6Ztawmdbg4Zotgqv4
T+SvIDslaaD/biMu/BtTchH60UmHQtgSAaNyIsLxuLRTuK0HyqVl2QhDELkG32CwsltpJvJ0iZHo
O/BQTNrmElEBQI0ynsfgVVLUynqbV3s5EonLZNjPXHDKh34eSrZo4NgSK7t6L0PoPskiNCj80wtn
HXjIHWTk1rNhgGvxMPZAs71WxcxS8D8nDvFGxBMxEEmsBjc/vLMmT0AdJjopAnF+VjY3XJ0uXTUy
bio1FAmUF+DvVdB0XXq9gxR+rkiAkoKaFuoB15Br42XHOS4J+mXyXHYhvQaOmrkQWHKdbe6mWzT+
gkh7ETRUhreIk0nh/MyZA82dkFSnjjXXNqgtGS4x0iCX1rGZFFBHUHpWmnxNwaerOfisrt2nCNkv
TVwJklex67wAridCTkePNniAhBwSOC21184J/Q4/SxhglaARq9Np6Sdm/PnxmiyUULv26iWYB6U0
OUOCYJ0nIIWS2oOawoPO+/vCBmP4qePqW/VAhsdUduKjntCUL7IhTp8L+IRh3jZCWP+a0Znlu9Nq
pRnMoxwk9RFLlNSe+1yg4G9w2dDcoNRHEs0WgDKshfjZEZEbdW0z2TJeqyeUn2f40rNpavAM5PgW
aTA+TJ9EsHoyUl6u1nGd6iL1v199ZSg4uI0DWSICFyVnNsnpDseEJUG9TkOIDk77PAWtb6JOb79b
XqvCdQp3Hv9j9oMWdr7KuiDGfPWJk2qGWXCXhJHkvGkxMsGcYuAnz9UYLzOgVNCELSUXUTKWEgYF
rvFhxQqQjU4kfbUk5OSxHxGIRlDyMpcxRZ3ZTPDWPepQDLU5ttkGMVEVKLk8lWafZV/zjgkvOy4q
smvO1/oHVNmJs2i2p+PDgriF5DUQdF+iLKO0KQhx2ym8kzIx6745TYb0fkwnbIy7qSnwOOz+4Zwe
KH5Fyw/6P+sLUBtlBY07po5oU+ObtbjmT+Nz7pOo45JLl7cEZoCp89v4Z1gLcLVD4od+O/8z058w
sHaTWU3paw/9qKfrrQoq/9SDKY3LBb6ljNsfmx08dloPIa1C6bCut1YVTYN7WluBySe9EIfKInlP
yeizkSSwE9yd5HfT1CH9d/hvKlKtV593JdCiobAKm8jmQvL2ZymvBGdegp/gp4xNJw8CizbwiIIF
f9yDx6NLT7iwW60tlx5bxzV713sKGHVnxiZZ6TkBqDCD9xgKeqIaZ1eLL6VHqlmlaklKTt6gUB3Y
7MG+93Uc7ilTRurnLcSCF4JdeecGKf3/i64NO50L8J14GrFGGCbr5P1DlDqWOWcrChBlTGdFnQ1x
P06leHPtVdUQjUvuF5ZdClGpcRBYdHPmp+3HjEKHKLNtAauqH1k6V2eT1ldcyAJ9nLUV1n0x7MrI
O+w3Ix9iJpnKb7HwALf/AsLQ1Zt08TySGCS15UI+iv7eQPndsNFiZcPegO/KiOwyhmxaGkPHuH7b
KS+oH5WTMAIcQRh1O4Id4e9botGTEKdEXrncyRyvGKismkPZ2CIUlLVTHn6ECJVvWH1c9BuH92qa
doiiCc1q6qxrT/Zj2+W6U5dvQhu7gM5y20ucl7Nlz83umUAdr1vjyFIddwei8rEKfxxOGAkfnujF
V85qUjoDtKkkYat7xUeFtGrs3KWlFxAL4FEaubzsCzjedEK7CWmy97FBKQDNNNoKXJYAuSgE/NOJ
5eMZ0NqZMmEZAxGgahq88FrVQ1HtxJqQ2siRwXNUKz6RSX34zVxTZv7QOxU+zpEhYN/gjRQjHDeB
n9YFsXxNOcXbACIEuXy3PBSjRMkxTXruubGJZ7alwPloupLtadlqIjBZ+oZke5OOAj4WhzjLe6Cs
U70CZdWv+FoTrUdAStAG8yPmirNKD5iQtnsySPft38NEnpxCpSyJaj2IHqQZmc9Xbf86rZOoF+6t
CWMttmhNwoJjG0liraoIZFU/J45w0DXPqjcKHjXJW6FL4exByUm0jepoXeTfZWoX/TqS8nq5WCCg
LU2QiEaUjYwwLGOJ57MUw2wh5bMZd9Of47WZVdxd+JqF7yknxIZm2JsKhJlMY51SyqWNJoPno+D5
HVgRAw5CZo9yT2blTbRca8AdRYBAbBk55bq7XpX6n5geYJFibR06n9kkw/2mFhwLzfuU3lcQfj+e
531WiBFfBcj8prc8cKYEniFrZmqpfDcyYty81Pn5QtJ5Y6mXCjVbQlVCU+AfqY0mjDjDimrew503
3gyJ4bBj6+1+t3qba5jk/vn1tcrLzTi6UgGrXtcot+2ok7sAXm7pZiY6IPLHaxxG30DdfDZIjFJk
rZ7kdx+rDpMVYlzOyrg52I0azw1tVTH0bJXmmotouYmSvEVmMweIZ0diri9YuemL7kYWRpasK8CK
IV3prIJ30YS4TOZfaHSUB5yeNpg2qsTY9dXtfrDWzDqjTOQMFl5z6vCKifnYZQ30fQjWXxUQrh54
sOnRnXGsoORNljE3J0W9glnQICV1OE1Gp8raD/8zf/tiRyCHlog36iV0yrck2Nf1V3DLQhlFSwJj
EoMV6UxUnPqEic3L3mA5ZQsFlw5L3Fb1N8JxyK6yHvpphBq1OH9aH1MZ+PXWBddcwTae24B8ewRN
xckAfueIJ5JXcgcqo3hfng7Y4ttgOp5odSVQHu7WylLKR4WOPw5pP2WRvKcTOZXoGVhaB1nfbO9R
JqO3RXlVTJbkfUcmzpScVb499JhmYd9NUiPNO6dTi51M1OKS7IXdRSRHMoMTp6PWQ6J2BK8DLKvG
4a6Kzum5Ie8Z4imZ00jtYO7TcsYz+yNBzw+1xyw0qH+jG6IZeTi/AyrVCgLpV6s7N6O0IkB+qrcB
mqKXzC8kdPKGV64d9nH8+CFikEXwzP4OVjeIGz5U6jvuVJcdNpUPYJT+Ad8HizqYUAB0nC3hoVPW
DnA5VS6SQ7hz5fZwVfWAU/NImAvI6TOrcnsiiedgV3vzxmy5BM/EAjS2FDSSef5huEYIvdwYma5C
UaNDKLcE7fslnd0HNaYLhsnV3vb4Wurk2OAgV1hQgghicYw6unPHHfpt0KmjQPNH6cAor5Ux0dSW
vUyRP4eHngsufPOpjjM+p9MpYUP9n/x1Ka0RUdEG2rX6C9QPAXti+R7K4gos/Jl5JEv1WFJ+gV3B
Yb5Stk35rHWt9OskGSlMzM0p6QFd+HKSJMMep0nvk+/soIRlp8SrRbmDCAswwrZVx6MJyG0LOeK0
zBhdyertG0/iuMZUSKcfGtXTXPb1dMhbiN4hBfmaKbcnt3Pn/4kSt+s+GMzArmzJaGSD+QtdDE1x
p0bcSrdJmRaEldg/vJE1X4CUhGRIBGAFwr9/t7eDNDIuQ3xS9ogk7HbA1so1Ugbhf4UThjhl+Ja4
3Od1fycLmjzP17FmOW4XdLO9Eu0Zc7MEtnQZVRLfer3tWnAK05fPEiEHIZVHS90q9+6tC8cRPly5
IeNtmMRiWVdeN6Ux9cQyc/s9/A3fn2DVIzvgTSnluApeW1Is4KQTONdAZadBmU3ZSI0jmY1N5buP
eAgtwaJKriaFKw6kj6Xq47UYjUEVDKRGqftt+jwi5Cze/wbpAxtEJyap/KufTVorRaf4un3VihZ7
LzqgITT6MYgNmetLMWZKTomRSc3udjRFMbKOAu96bKHuBcz6kQTfHeatboNX5en+HNZBlf6BJH5z
fnYxvZluODwzAm6cnHAfOI0TPxB3P/BF0PSxYgMuJQsCI4xijlnMC+m8AnuImo34Oip3fB7NCngv
+yLQ7pO2WWW5gWgXhtfJKl7Vz+k1vo0HYgnpZt4To0oGRd74UY1gPzAF+UtNNxuprPMqsEEeE5DM
i6p2N8AaKZNGFhNS01BwkOJVgrpOYocwJrDrEcjxwsY2/eGVONm8SNk99e8KsHE5DwVhEEV5fGH7
X4pZLRfkeeIMNFolCpSExOE4MuH3wMY59V3w6cFWd4/GaLXdi4QptVLdxCZQOwxP6kCqfXCFmEJn
3GdSDj3QUTiDa28+mDA+S0Ohwi4jVb/KU8Eppufgt23Nf9DJgtYpeczId1aXMa7r/s4QtBUKseeM
cNgRsQYu6CJaJFYFjaaILp65WbmU3Lg9utGfq82r1tm0KmkGIPh6Xr9SI0fAt+cbgbumbaSZGwlK
y5NDuNNI7CTQTESda1VASJ3+i2XmAAgafXnVpDRSz63fO2Am6Oal/wGQjthcBNlljzZafCykGeO9
I2w1N/UBnB5FD7nlhFNb0m0XrcnuZCUezpP8oOgnkqqIgD5xmmU73oszfZ6ISXau+9uuDGZf43OW
AJt3KQAmlpFvs340of/TXHPgPDzpsHo7aNCsdlqDwKbY+4CZc2tTnQgQOPTpF5oVFNRwnz4tVV9I
IwZ7ejqhaRCbSWzz8TdypLGciTdW8IAcrIhEOSa+CGF9MYfgZO1GKyswrBA7fpIdFB6iARwwwhu/
SEmKeD5IXeYg8NhbtbFzgVscsWf5djIVcptX5A7tIgDEgAZy51HGxhs3XNYgMK73BECRDNaDdKHS
ynGjiW965piJUmaHiFVzMucMhd6+L7Sl1CaegGj2yt1jpLisk0sRfdgt78yHrrA1TntuHTpyUQpr
oDGr9+hhr9eCpvHvVUgW0oRB1wKf9+JOn7jocVzHjXQZyB+zJk2dyb2pL8L0h5h8d8JVeMJ7AoCT
XcqkmbsdoWgke8yR0/1BlCDnbj6Lk23gkEO/MaBwGTwiUV/ZS1lpEUqAcZJ6FXFI8Tjxl5lmmIxK
vog9iB7tq62dYKfH5r+oVa0tyRapPgR70xBTQmKLDy3wpUzgSHuwuZyuoR5gbu+kIdNp9ckazU4S
KyuL9CZecMUpJjjhNwALl9093hrG+onhcI+TRjZgmkjhv7b5DuHsFEPnkKX8L8VCHK6TeuARSygy
svnkav5yB/4PgyRt+XJNP24NI9Ly5ISbWn7lGIClpfFMKh18+lFZ5C8q+uvFA5uDoEmhPziugXYD
TWlAsC5JzdLHjCwfxnDrTbJt6j8dsVEpK7jaMYmfXQvCFnaleBP9irYFJ1cu3UGa0UrxE/ZDk9SZ
AmKl3IK142fpiK1RhiFTHC/pIf/jPLxhgHaNLvasxe+H2k0FBcnbOo8TeZX0OrkGCahzG6GyUXxJ
/G5nA6lX/pQVkEJl1hDpLJYUo8tobn2cf6wrjoGYzzVpaB5wlcNADDSiPP45/410HnXS8n+zvvwT
106xN+8bWMVUAHnWg5xmSYQHAZuvjF/3zdHB786XDMI7FEMrs0wYHXkopGekuGQ+rr8YKZeK6bG/
voW7+lbFd4Bk4elhgQftj5j7gDelA5b+Z1FMTvRvuLe86FNAsFYSL0Ul/e0O9jy4OTPt/93ii0Y8
qvaTH7TDDj/mAxyu4GRs2x94Y1tS0eXbwK5qiY5iF1L+SM+HHUIsmsM0v9sW7u/gmC+lwe8Eo4HX
2oLMVHpbWdp142AWv0Jy612jfLBL3qUxdXWDuqNsjk166at1AHpfhmn/d+qkKv3Q8j2KBhtJ0M3c
KmduuOWJK4PV4+sxbkYUSvKHz2OUinKdFIRyIvs+R5Bwis4XPrD/jQ7j8bNYXxaVGuELo/rIHqj9
cPV4Jx/rU3vtQurCTcEvDyxBU0IK+dQnxOOSZlFqPpsHYvcOHkuM61cqOvwjMiDaD8N/O6cnx2w9
7CbdsQLJJDpD+9bgI5CAlwfaK9Npqvv+9WmR0DR/9mrooAdPpNvSmAbHXZQicpRAFVyr8HHhgKVj
nyv0mLqVqqJ+j3WZ4kcdkIVT/BLK2ETEwPerttNo9tRxDpK1DiEfVf/jhatuwW4WRsDz4kp9dYLK
/bz2tCcc4kCNmkFFbMbfKduQmyHGAAtcebJzYHFej09wdG0CQaPdRmdgUDCjpz1lWSj1PLG9kVfl
vjrAvpssppCAztaPF7etG30JwZozXtSGVOT5AxPXi479FP3JNsc3vOxZuWOJFPQ7sniITCjIVz6m
m1f+LygMboo3352lWIMk9g2uzTzkP1bq9Lki5GY+ygUvRGzVfJHDB21tWTNFeh2Zb6eziyei1iDp
822iFSDUPiIxh9sc/D4ILmFgrrg8JeZPF8j43X0vF3ssp9kPfbFldZiknyMyKmHM65YcW+3y67W3
RZX2TduTfSKFA4Naoaezm5CcY8HVzmt8NNKdt58e4/5Skwf0fgcV1aSegUhheEU0B0LxWmSD3q9n
Ly8AVZyca4t0h/g4v82eAqzGWqZjDm5y1WhqP4zf/5bdi3s6+SHJ18wHEWrXk6u1Bp6O5i5RC0A6
bsSkLFn2IKu1/+7RxrrksrVtO0YsEYjZEvMAyS+eO1qUIZYoy2y12SyQOoUFQ9/bXRwJQlzBs8iG
o64faRIMQoOuOLAWPAhV54PVuioyi8ZfkcWR8E1QBvcLOvWCaUJDlpCYF0Fd43eLq9JUduytUivS
bJlcjnNvHPDE0Se5UfsHb3/gLbflZFcd4cFMIj3IDn9uqS4G76PPiGSzlYPKMIbvlvn6+qVeWmFd
FALEKj6wU+e4NhuAHS5bs/QJ1IfOd2NkiL4BDoljdkRUW9r/7EqKoR0qam7rhaON/t7DJIZaJ5b5
MekmAHTYCA19n/IEd0wdSvK5dmXLk+ZS7cjcUWQub24Gy110+y684rlD1Bj4+TMKeYVcdbrJBFkb
zkmssKt9jyWv6uiYAbAPRiyRGvEeki2zqTdZk7x40x0b7bgULkMu5qoPoW33z4xOrslYF9woxjH3
iZoek1aAAKY76gOco0GbBm2j26DbAZpHPoF26fYX2P8H8o7n6Hn15VzWlaOlmRgVFoMT/Wd+b2tH
SS33R4x6YYYs1bqevdbOEN0EUCJtdEaVoBHYjtK1jPCfdxatn+DoGjZgpyiNEdJJUJXYTouTBmoI
w2JUlKakDwX3xeB6nKyTRMjbCGo/XCrCeilalkY7LBpva3Y5OtT8uXs/eyv15CNbe81eZlaLXOiX
TOaVDGrwY+OjRNbGKRc3x9iZEVZIdvodkUp8ehFbVhtgjcR+iPaL1lHWZeggEteROWSHribVq5Gm
pH8Ov997BCMdTGPykdH/c8aCTZfz5ymB3g9SkJiyAdkr4quWpZZcE20d5Tx3gDEtJePmEHHcsy88
zdg6j4OqZqOQ58BlRRMUAcpI6cra7L4SLswB8a/6sKz4aKfSNlGbGGwIrDiV/3yfX4AZPkqoGwi0
585kLu4CMn+hOWRQg/9kjkiPpx/hKx5sUG9slQuYPOCBHfD+hi/vpP/EhguPOPkRxv34lRf9RhCc
7adb2I8mfZqNiHCLNRv7ygynSVOnov0+ZoxvpsM1g8Kf9vDa8tWgLN+zmb3P3YtIPp5+Okqv2aDC
6GzW3glfJ9OrOqD4K2/m8UUltynL2xR3+Kpxrin+HTIo9Xr3rrEbYapFiPdJ7ngD/zckea7ZbN/E
sWkBaO+twHJrbjKOXVWMn3RrF9FNXPnUBS9rycV0fM59KU3PXtRRpATMHXXTyanq8HLpimikR/zB
QoJ2uLdw/SWJh8zevkpBFhPtkBaetjVACKBas/hqmTbeK90Ab49fchL+7sOgg4pem2u5wryYu0d8
oeQuYB8uF3cXed82cfB4XC5p4U5XfH8bBTwWAP+6fI0zsKLcAj0FOy2QCDiustypl8ratmOf/+Xr
rgsSX733qUYrBYp0VovWHq/FJ9qhoKvOOGVKw8vrGkKAKNF4huNb3Km38Bcu1+gKItsj+xtunLOo
8kmtsyvW3dcF4bH4kWS+X/XLVrtx32py/8FjwZA3p1Kb84quwR9k4OUeI4eO7GdXnquLpgL1p7QF
PdugXDtmHcdSaZBAHPX/WksmxSONETUByhV94VG5Q3bnLFGC0JNuhGnNIFIy9KaYOonyTtnffyNK
cvpiKEoBShq5jCHUDI3aL/KsUkxC8wP3msclFQmqTziEwS5bY5ToKVbX9AW/aDTgj9VkQ29Qf4st
JCCtuQiF0t27Ed9qsl2RcS+94RQvTkO3sgomv2nBbnA+zioCMqt8zbLp89c5PGrnsMspKA4HlZ8o
lb6/lYjNOSb0s4Kz+VPBX8p6YOyj+Tka6Qie3hyvgkAVd4PKD7zo8OiECL4AMJr8Ev7FwYcq9Tl2
PdzFeSiy3B7Hodc1vANqTfzR5FF87comRixUNFjrt8/ixauyWmVtxRmcJEH6quUuZEUwVV/Hd8mJ
yV/946UH49XqCkulDA2dcNCpaI4N2fTS8YaXyX5qs5jdc4pMh7jI38V43+mBi7zjpVXxeW89h9KA
7VlRDb+9t7AZy0xDCUSg114LxsGs6AoRA5BhFUmdv68j1Bt5Qersfdi87uWRR1VnFYrgMra6O3gh
gdNT+WeSQ+SWaDEZVcm5KJnK0cBrbigAOWP8/2og1Wi4Iqz9ZXmdVDJfFVC5Z+aHqqfMrVkbRKUi
Cn9nQqW2/opbNITdfDYbaRiaTK0ApPGWaerl+rovP8wmUkqE7tAwmpfVlhWONE3PW6Rq+6YtvuzW
QoUN7wzU70ti+36b07uTmUTDF85x3Y3mdAe01/iyhfU2vr1z0JHbPn+Zgsxa4FWIYCskxBBkuyDd
D0KDWaKlphdig7MeqExE8xLumP6iYgu6B3WUEBf9QHX3Gm6U3s7Xkjj8YMxxXCPuNCgZV6QyscWv
K+hvR9lSAxYJbUulfLi5FwWQEaNq4+2Rxk4I/RlOE5F2o2LbrB3tqZLvw+WzVkraA1irdRGZeXm9
PkLUen+4nz324GkQO36B4qfIKeYr3w6tkN8jDVW42Zqi11UmNWsKfVvJW7ymm7feU1AAibtumf1K
ot4hqhUmpuxQH0KEBpYVYnRrF4Oq4+L5BReZavY5rKdyxkdMPEZHoYiHTur4F+0hnGaWT0sJjcKy
74Pr12j0j9qH8AAHouhKjUj3I5UUVBZTX1q4TM2dtbcW3DsE1/kafxnP9Wfv0QMgJjMK3VMUNrP4
XkEJ3KB6HsPqSE8fp2iT0qqL1n03IGyazGRFOI1Xj81BZmEf4KgVdJkO+NDHI+8HtubYOwYaR9Hj
U8qr+OPsWlfEvo7b+9sTeTPzjYpDE2XqD8JxL67+feC0pK/lgCENe0esj0URK+mjpHxvEJ2kCgqz
VDd3vw9nH2LCrO4QEDeOdnXD7gojxz+vDtGYCZZsZlXF+32bq3YBC2wZzC4T9BYh8izir1S4ytrq
Bt5B57ngchYXbDZQTJqdYYL85HEF4qA5DGywxWyo4SDmUi093wHbyVfP2IYpxpK/Xqx/lwbviybd
YM8Lj24h3Dx22Jw15SM0XwMl2imOpFtoNm+laYhZXDN0c3luA+nDVydsl2i78ujcrDkGA9WzxsnW
w98a+kWmLbv8Tmjd1b0rewpTUtnZmlOWrxW4L5LbHFqPzkLWwf9HSgNBFSF5DhYdGruFHpY1XW/m
ZAYhPAiXC4Z7EknnQlNy6quDFOGpb5sh4/jQ40pfIqnCtgH/un0W/oNV4S6LJoY9j7mTC9F+VJ3T
Jk5cW4/DxgY/QN7uzJsPBOiSHC4SBEs0FxXqe2dWUvv2BvTamcIZoxxfC/GlIoo31ELbTz+CnbdH
9D8IPx/NHaFh8ujyksNc0J6v6qsnhkG2IrICznI5j0edNWFAU5X4uiRs0WlJ1HGxQWkFKRIJvxCJ
H5l/TmqpV2OVlrl/mqqKuH17q2IXs0ONKoaC794haOBVI6nc5adBYgG+rIbhjOIjghzaq6XFykRz
1RiWzVWktWSdmIZ6PRnbXhAVSPfcT8yli63NYRZjpA8Hld0sRZZJaTg4aTfq/iWeDDepwK/FhYXx
rh0MhUqIhF/7hsABujspFQWnHMI6ap8KDRglRIhrbaPx42wrAHI2lNij8rvrHGLBlqOTVjiFYqzX
I/xJRXGsnN1R1LCbLtrqBb1WqBNTmdHQbz957jpIyuxolUVdU35zsdvW/zeY1XH92+sIaTVOyxSW
7B0Y2g04Gegsshh6MpCtUaCJjni+/d+o8a/hjsxVVk9fmBq+Ctc0P3dDo8FDcO/Enq1XJVd5jNMY
dkuKYX0b1XiAHzO3MWTSxfmrZNyBrsOBHMSRh1MP5BZ7PE+x6yq6qWcJr99qvS3XJyZHiAclNdv5
pYnQj2XwuiqKdRDjKMpaHSNweW3E/+5WjPC/UMOXs2iq3SAZiThuT0QhrTpqmUeUWfZhY/tPTtMC
qDz19QX2RB2ClBYYwnrUlZjRl447bAyoANINgvu5pjMdVkMunsRoNf0M5hTS+d70ZrYALJx3vMa+
b3FeFzYFVmLGOef8XOgQqi5z71TuxhyFcyHb7C17SV14syfI0XcbsLay74uxHONuYdvAa+L+B06O
/RqBCDXyGMuedtK7SqozrpzReamU8X/le2RXOb6icm029tzl6MB9y+qcKQMwtjisSfAYNwPIy/Za
YDto2+ZZG8+CR6ARqi6cvgO2VxSG4iz2G2nAdv264ZEeBccXtTB+/CzBALiwHK7357JsoS1Doyan
Q/+BToGbvssyiMCLgSeGlsjRzLU5QJj82toQglRTGH361ENdhZLhyPN/XWcIcB9Jo2nsYlL01qxr
o5P+4ScMa1bniwcmQFi9R14t+gCj3wZlfWndVCBIbUvF6cKYDVM+S3L8UBXHetLkhYjmXbXrOkvG
/aS3sO4ETYC67PyqTNFSzKwFGI0uWTm8YbXr0aJ31TKerJClWtjNmwmXhjSOoQLyBK5Vt2v1/ulC
ch5AAmqgCC46/dBB6+PKl8AQM8BbOsWyMGNrCQLBVAIvdLWpb3U7a5tfLAPxE5LksnwsrqWIwMoY
LrBkOBsLzpBRe0vKZLHBloYj2QlR3dlTbSEDriLYVF9cZyEtwW+0LvVsUeHAiY4WGxgBrzokGG60
Quh0FmAtkh7Q1IuTWRXQ8T17/saA+20X+UuZVgVtjI2aoknRNY48JNW8D0/XhgLAHS3Sp8L7BwN/
iSL9rO4QGfDn3oZ4TT0WCBXgMYy+hHPhTkSMjXENC5hKcTKJyOvdEcPefGg7TCHLjat9JNYV9uUW
ZgLJbAMwRrJvYQrz3OLEaexJH19J0RkP0XxNX1xxVhi9NC5oMXzQhzKVMqKzCYY2cvOx7qGYTm3V
8lYvS3Stw2+8nxdvXQzV3p7aLGAbbtxi8utHlM8smDHnHLI6YfNLGiXgRSkeRgqP67xXHfqInl58
VCid/bPVCA/U65a0cBeIgqkvqA6w2K8MWWRUiKf9H2YZ+QxDk/0NjD7mUqZ7sXfZa6Kz4gc/TQZq
STNIas4WxoDt6CCeeMt3Mhiukp21MHGwVV/4n0y14jWh+66xXyYQKr9TXTL6/A7mZkj+pnv84JSH
1rK++uuhP+mchurT1omXq+JjZv0cU1Qd8SjNz/vBIzwihjwfDPEx8uHIsDODsBfB1leFA1ibct9A
ctNmjtQZ8hsPxpilh2tcA1ifFwyn4rd62E1innC4Sdq8c9m+rXp6XADVraey7bK0CBEfldFSQeZH
Hxan0yVBFts0kbEeb32oKcGcBxKffkrqG+FX2RQNF7ehpoyNQGfHS8kRfRhLSxMCqbSP70hvs8Va
heCyTc4vmSZE6kKYABbPe8WI56RZrDZhRfPNxxlZguy20Ytu2lfrr3fmtKQtZTJcx4LvTwBog8O7
Vujc0ijnpc7DvfqHkj9wYb0ABvGsbFbettjT1pXF/wmmlTFvWUFDxcFyaYaitM4XP1ML/fNNKSfV
btM65XWdCNklOHuDwszSvnTW22/PYlHeaoigelC1u6f/T5ZwetD9gwQU5KFD0R5xvp1irowz0VFd
wjErIit39n4+hDOpLCj4vN9N3Hoy9NYnOkLwv3jx75bkyRFM+Ht1/zFNcnYeDkfPraVmt+J65+cq
r6IfiR5+vDLdQgL8OyFYZNAxJPduaNyIM4f/SgJZYYd0i3RLJsiY/NjYbvTRyWeYwuVn7NN3ZkBA
pQ+usbzH3WVoitSzBASHkh6c4YdPa0m6zzzKFTip3ZWD+EBwPrh1LeXisBoRzsah/iPGMSXmpPDH
MOSKoVvj7xoQG4/I2SWjLEuanuqKnq5PMENrCsUpUiu/Ir5Py9jSlNPXLCS8S+GwpCYxc8JE13IN
g58b6daVWxlYGcQ3AcouiruxiGDzPYUv9JeNqnIKxR5zGlCyA0AzB2O6JlGj37Oj+DgqHCpu4+4y
hcNEl6gjcNwRCVIg6P1JneC2wRNVgUs+v0qKejsJ69RP1BvGXggOQdjw3CxJI6LRs2M+wv/LjZhF
xYivIoLfYP5nvIkUePO1FaWiFCa60XGlvnBaLEh2yWbyXCn4XcIuYNwGvqHlrv+xraDiTqk1CQog
+e9cdgR2whg/kASBW1RDfJP+MQ+5nGAP4O+kQnev/HWSsvOWkoLrinbPxivMN4R0rgFmqaYd44hn
fvcFN6sXnRpmNnqSogSt1wQeodUBSagAmwqcVWSG8Mfp6LtGUuV2suTEnj+gVlg8rQCHwsgCBI8S
9xzzgapji2dfEFKStfVQCGlojDDdUei0iU+rt4WyxkDTd3Wz4GzRonP3UygpdSUhsORysnbJcrkG
j8CYLtCG0JhScHIirttnNJ7/tMB7eOkPuWEnLGUV2fxEqfVWOvC7SeT0VeJLId9FeyBaI20M6J7L
2C0Dc5MKfn3vOvEU1w5vsAHn8nQLP+6Zqtg6ei2EVFPKOyol+OMvJzCgZk09VOtgA2fIe107Z9ND
gkHXgWnFfCx7rAmMf6aoWBbX1iNRp24gqSnn7mMvO8IRFe4B5Ufv1QB3h+3XcDiB9NBjsls/znLs
Ewm+tGeSSsm3vG3q/oHNeRp3I5At6d8VrIRyFoa/cYPAZntyUgST1QioiU4Um/dk6Fbb93eQtkkx
IxZJA93RJiUXOVhm7fcbpp5hRQfGvXmE/9dx1v/E+l3oL1h2qK1abN+3PiZl3Y5IYmRILDxQUFD4
Uq8J+c1w/q5KVuRXLiirxfClP/m0LcYYCrA6wFNQPM7bB0aDzbzopYZBBa7wkYk0kvS/LgK9Pjwc
V3SXDSRUmAb2R+iLuonnlurQnTtfcyAjHNZ18E9sWpBxBQG8TmrPGOXbwKBpdaBCRHy+NRFoojMX
0e39SlVgtyC5QOtf1kh8A0N9ygSO4wTulS9kWfGP5L5d9AznXKNqKwqSOnAsze1NV5++ByvhgH75
YeZaT0uPf8lLlS1onTnBoCyxxlfdWYNcuhsNA+kbH0LIyA8XeM8XCDqv0iVAZuXCwaagXsgTipnm
nKonEJ3qUbOtnGUmFiGpjpsb6/pUB/Oe06bc88dS/8/SwW6pJ4qj86X6Ll5KWyIPRRVvQHwpHoOJ
MH5gxs0DDgeJJ6s8ucZiqvwXGGLcHecEr9aRehsoMIypkwc72pLxr9HjBNFGalgY5eWEcrKBMHMO
x95/IU0M0p+LhW1sNIWcWE7TurEN5nlz8n3p4ZKw21upGWgAnWT5NgCjDeZzKn1OpudwqqWp7RvW
eUtfHI5oE/ylgXjZd/7xKyZASudwn+Bnw98CVkppfiikruDTCof6GMbzEsi1jEpDhBuHg5BoOZnN
AdBbSNeJ6bYEmBGlKYxd0ynxjpuWD0fEx+TtphiRGge+OAs/6OebZLNHdDD3aSoiBO1JCRdHo/1W
IB+ljtFxbYcEimiTHLhZ14gIHi7AyLbY8aHl9Vimfa5VER7MwvfbEHfqv4K9QPlQ4EspWLED5QNT
u18kWDoPhfOTS2mwU+8FwXcYqfRy31KFHrdPgcQezh3pmVizjaLRDWHeRXZ+0t1UkohX3lUM/OqW
K0ECqxMm8ezqJ0jdcYKSOB7TtA6rdBvoGOgDPM9NDVAL44a/vZQ6odI7rMzd5WAFZSwfV5/n5obt
Rq/OMaB2GL0fupZeNTvRBqXFEDgfiFS7L9tGSLF7iDyjmbGVcNK6KPk9ex4fce7OqZmOLwnjwwiO
iFbNk3ceVtlf4twQhICx8bJhX5OR9sCumVR/68gd1sHgSEfu6hn00XDboaQqlRtgIWnJ08pbHcKU
gCDT62s9W5EgL5hnlWIVJeEV+U+r7RDIVQBAHj7x7iMgGylBjQEcGYncxrkMV7FQhEukH7hI9NRF
kd4oicClRlt/FjdJIX80gAhxNf2Y9BTtdJ2vs0qHWhya8MkmYmyKRqO6Z9AFQPPQUuG6SCstYJBJ
f/e+DpIe7ZhToeVL7ZEVVgsLsNUdz90IALvY/hAo9O7z9Lsmdz9VVR2sNbcAZmH5iRlxOVakQUGI
T/mXvdhn24M6LQJgoHPFwBcWih1sJuKwuPjF90B2uulvQF8dkKRiKUJ4oX8Dn4yXEeGchvcLyWcM
ZSceK2UMeOo2NAvjJTV5vp5Tf2oGl+GnNAuT8+ART+pAPEDQfZyOsbzxh0eGzAdrgn4APurrhUhm
nA5SdvG+KpUQ8tA1uRiVZ0fxa1XpvDctWKNWzH5YATxhAa5dgzXTxwkLuA1IpNt37DK7E/BAL6Uf
cILSpxuSQph8CXDfoJBn8n9VQ1pp7riHlEXfrDDaqw9G+zLvWZKuD3RIVwOWxMTA+y06uxU5vd9q
bbiOuHjWm5rIAT1pY6iYCXp0oasB7u/lCVE/wq/XNe81SHD74fbgUhNkseymd1nnJHJ3Qq/k4ozG
bdXB42BEMfaW4l2H8N0YoBtwliQhjsDPabEx/ps0iiYp6eBhTO+wP6PdovGxNEC5uHDaVnb5Z109
Dxla7pbyLEoRRS6mav+d5AyW3DKOwEraKHSMMjMIqM8ld7U41lPA3RGlsIapFGOhkeATYou0QshI
TfSWwfGFkP/B9klDuF3rJW8TXXQ9sCTcOHf76NG4lrqf8YXzjslpddP7wQz6+hARGyZzNXZpoUR7
fj3gDvHD6M91M+9RgGQ20fyzzZj2kruG+wCaU5ZkMjraRbdH4qupIa6OyxTKZJweDCIbK4C7Cnji
IAdXd46Nmzz59AcX2ac6L6icTS9dQfY8S/Kvq3Ia2haZOHcrJmMtyTKS8VWRtx5yUJbbkVzBxdKQ
8/ard05wTn9rcXPE0A++BGeH+ITbq3NekW6Y1qiqvf12Gsbz1ddB2onaPUtZgeNva7ikIuWaa/2Q
TbouLy6WZAepSwDttQx8wavaLrtLvCcvsdqMmHFwqntrA3YmSznUBBqZi6MzqVuxzqKfhSmcptqy
PqZn3buA8YmKgFR3nrenSRKdl+wZsP8IK4HBPF1elYHUwu7bAAD0r5rICZ3G2ax2Bwl6U4dKRTRf
yEhl/fimM5UUyi5eZX+wzKeU8o0kCyLWcbn1gdrqvhx8xqC0ZQdQ/2hX4TazZ9s6s2kDKl+FrlAO
7jrNTapHe1k1KWEKphjB3CCrA9uOTWOzySHzXDDUUfs9pGmHJwCI1yltikqkaAUDTU6SbYa8BFi7
+zpxKMu1bbpCkiQyUM9M8sDSln2fr2CDF+kwgWHsI7FkB5L0GLKwdLCLLPaWeYpy8lou4tgigELM
tFFQzTXwFrWoHzQeYtwYM+HEBLBG9oEA+laRbVI0xK5vIZVI0LtuFcEaAcbBp8Ly45L/u7cx7qJ0
RwwahX1bO7H1sNay4kU23+ueAZ4TmjT/FX5zc+HyUtsjzpvwg/o7gf5urnL+MSvhZc8Ydn+oM3AQ
Ckn+PxE5VWmI2zhxM+pguHD5GZHuep+zWlN2cIWdewt2TC2m8gPZNUujmQ6w/Pwe3bRsrLs6g0Ia
kPwicNTgF5OFKexaUuyJ9Icu+4M6NWdVaI4AinaDY3bMlQ41jyQ2f6PYiyrrA5ZHKInI9EwGT0Xu
JT/qFGjfFxX8Lxd3zpRLydU1nnuTqugaK3d3Jht9bZUbT+oYCvS0n3xenxzNJyso3krsKrfeHW4Y
YGgQnGIXjTRtqDfGV/I3aa1T/GCipAH3OegvpQ4rDAu50Zcg5BNmQjEPfBNnKUTjICpG3IUZFH2G
YQbSLzH73+jCXTQwadI3LA5wP7ZM4zgKLPd8jLS/AWrd4+BQ/cTmnyooQCtE5zqDnNKk7ljuFu8k
Fxoukk25zTrRR4AlpgaVxlSoO69YsPc4f8g4nHXAB3+6fqW7hcx4JA96iF0iRh7w34vqaNB1hJ7K
NoITlF/E38YGUNy7wxaNNxGzVEaKqfZ3TMUr2gM6j2a6tMYsZ/piyajcNFLOod/DhdajmX8xarNP
6vbAtwDK2soU/tO+9Z30Q4jb1p7TQk2AkZD0Y7PVYModZnvA4Dpl8v/R2nkSslMIRRQywX7m0quA
FHhK8CVgP9+Foi3JgJb9OSwqMyynd+p2hY/a3FfG+12OyRXnRgopmpyiEueYyoTC7arqi9SO6Lbv
QiRIbTdDfg1aetOB+15Kumrrqjl91k4WOmtcHUTwC47ZiaiD5b79VNTUsYBGcoFic+BNHi8d8c5g
pz6imMHkD4yQrN8wdacwYgMavFKOz8ZTcz9WNVhNnv5ABQMqeZawSiEvimFT+A9A8367aHgMUNNg
Wh0kG/juJCfCefCl88dbbvIdSoJhHIy9MvUhAmLGC3soXrnfwV0KBRHFcl//4h51sG9T5VB7KvkL
SVCZPuJlF+ePzJP/bnffqGTgFIAJha/2iJWf6fJtxyaeQwsaBpHmKQaQRsfNGH7sJy6nh7LiJCJQ
aAzWf2pswf0BfyWslYdjCu1K85VJoTvXxnRX9Da/6maexCm1CHOnoogERjcQDNOOuUfHWU1Tm+Mk
Lu4jfta20m+RucgEFN9jAlFdoYUgFZbP/dLj3h4UFvaso/A4T8i/6TxbU9K/VB3+QzVCAm9O2QZp
9iEhmyL8jTcldwsQPO0rV27U/HtFUqwzO7tDdlnMgnkopn9Z6NFobCSFV8e4T4og/SulSOCoxuiU
5y6CPfzBnTtqQEuNfzpJ+ZeoInOYb52SNwd7OE4fJczsYMdKmXHv/aZQMiIQM84yphbM5Di7sQgV
sLLjRNfHCrAP0X9EdndA6cNc0eshgZwLoD3HbD57GlTYyNmO9jYnEu2esZbMF3RtDggFWOdHr0h8
k/7zX+rIyQfZsK3AdqttjWH1A/7GMMPmk9CgXkOADW0uy41sHIBGDnPxPAqtBpDxmw0A3X4IX+Nl
KPZsJmHMceOllQ6LAtXXqau5Xsxu0Z26c4THRozrej7lhIlngVYJWTSc0GDyIzqQ/T91cRwhVOzF
jQu1vNSGCs7JwabWJakZ6hx/k59699yqGwDJPof48FQjb/1iDvCMZLfakrl81MSQD9GuGSdQ+j8w
HJ9/dUV0eSxJubtQeoOmfzeyYcsm5j0GD2KGvQ8ccXM/IVv7SFrzboC/RvbnkVlCfYDdqyIYW/FG
xBaRJY8edpfvhB3rjM8NTe7dF3HEnEoOs7HZvXBxnj9KR/r6b4oqgabRCpGQB1/U7DQ5cLXviZnI
Ig4PzQk2bUQi098mdOoiVcoV/xAyh1cGhG6HUiLPTRfrm7Lz3rXTvl+PP4OwTuklCmMBg0j/8WjY
Pi8ZqGJEXOR/NXtRyPv9mtYuooaaSxxtQRANGqWcZrBpoSCZmhL7p6xxZGr26R8EIC96Oy+3ddFH
ffNDWPxdzRmi//RPWalyVdCsAmUX9DlwXUKkug6qmuRfP49oLAUV0hrITPLcj9Jq0NXiuAP1QNY8
WN17ohYQdxYlI0labjcRx7KQAFizrL+dMol2HoeeXHBJeNhHbgLvEUlF8iVtUw/9n+LYg5ZUyUya
cXDwfBwrZx+axBYL5L7kzVWpDk/qGMnLGEajCupdZkpxoZFkVgHUXcSlAO+Fq/CWBe4R01ghAYN1
ieLvDB1vNhd52J/hzcLU3cHg+sNSZyiCRge8M0EjVu125f6rkF7Kr6DqY2VenSKiuNGytenKOhzj
iJaMspviDq0krBHEYfXTC0B5Y95dA1SHZMTQSOlrKQa6l8TpTH+kXqrCrIc6y3SjmK7X9tGUmJjj
g0GzZCAlRzJYu1PuyB966eCGwOb85cmRHr3JuqbnWGgloh5yhgBuQdVXEeSKtE6b2Zbf7UjkeuDu
oIabp31vgcGr4mgUqpLkJbSg+HGvgsRrPgRHQPM6AaBRhnOrOwax/MuJmovAMmTg9lk+N/6Ififw
/08jqPMOi730WCCenrGpLmEi2vSFS9dipoWiyO5Cney+zLPVqogBlIms0/6R9fzKy4V2R1WWh4v4
DOyVRIU33+61FkvJcvFDMRxi2XOvNFPh58XWx64t07F3LFli/qCuiWgbrD3Rto+lFx0DrnNHDyN5
E4r9n8W34k42aZHSZMZHVYXKkBCwsbj8MDnoRaTo1XXZPgMO5ybOp74F0HqSf3OldANMM/l9OcPc
A7A1cLeCpvRTyc+oxKgfdFIIXYN9O+t67JpxawwMy+yxEPj1pSMIoGWrjOWQkr24yx443Hl2Vc2s
yrZjGzbOAU8wyrkeDJG4mY+19j+ujLgReK3dqM3FsfXdVOa7yOswFLlMJNtUcQ5oRttXSGwDAX26
Sn4HrL0V+3/AeBXoaROnchSfYZThnzO47RoVdR2FgjMmAXNaBcq43svAwJebl3FDdPxsXBVDezhX
BXJ2BvCSyCsexKa6walYovLc6K/7DDLk1hZpJHUAkpJrNNUXoQ8ejlb0PZs7VEMvci3iZRKEAxmV
Lec9b3JnTjDvYtPU5Im9toIZQq+bzKw5DFm2Aq1knVM3MIbR8Dewxul1JSyx4RWo9dwXTwYqGZLS
kPN/J5ZfHhiNF0aQYBN7JzoJsnIiRhacELma4qbIoGMZo6kZoteBMbcMfz37U9fZu+86/u1mgnWi
m9wrRNhOiMN4+s8n6xAi43uKerVXP7Tw7hDvdEK8/y/wzdmvbKozt5Gk8zMNxfpH/Bgisjk88wLP
M7+azWSw/i5ppQE6lt53x9ZSGqpMvesVWcshtbxOZ7km1KWJwFL/FI9ifU/5Zjx/4BbRQa9vaFBt
9iEWIpko4SG3gEaDPHl2twXIsSmxQL8MBFlsNICvrJPTtuO219xORFFec4fe+a6AI5bnKRElZ7QT
FggKKeu1BbGNc2EmmTcNarSuFdlDrz0RE54FZEtQwv/BvlPGux8pPmOWwq2FdFoDQbcZal61qma/
Wslq1enkd2PqB4pyHFAxziS79vwE0TKmdsF3IpvNJS/22eFY0X7a/0oDwh3Dg2GVKbPR4SIMWGMW
Av5mvdNEHoim0NJAAA+fhz8YVO1wVh5Cm9zhAj5EfFnFDOKyrSvTrdH/vR9b29fThpHTGG3xd8X9
c9SDelMSs/D9wYPglreAdcJWm/FEkrxKRJFg58mTl5/DeyyW/HlKjAmBZHZIEriv8n4hrZCppR/I
lN3ALnHMebziIZIrg7bRv/eQDiOPHC7PzrxGw1EpBt4oxmjbqjYK/ClUrvksm2yRJpyTDcoAp+oL
a54NrMMZtbTktjBe/hlyrKLnFqzfknx8HzrFgqq5wPjXDmUvtWtC1u2kGgZr8OrNBRyOLUkpEq5d
s657RYp+Vk12KXAYdTxQ5bhkP5DtYAxUAjazLJQujW3xu2ML4FUZtRqKHzfasZ6Hb++gGgUzPZm+
NlwG+2Ljteg1x48MZJR6/LtaptKPpgZe+F5Nlcxl0aO97oxGf2YHnqeakVHbehztOUC/jVcGSYkA
tBYQX9YXKyl5OIf8P7sxf7QzTQbGO7gtXudd1GJSXd2Vg7zBY6FXjhWtFcOdMkG+qQCE6Y88YzLX
YZ01OqI1g4dhwxdKa38wFS7ihjRZqFbq8tzuxJjeAwkVheKIGopVApJGxkZKVV/XmNtgaGNTIDcT
By9WZuc2yaKsYaqnkzqlXxIEadmc2ZSNGJDej/b8VgMEDbTKwehtfCuSd9wtETvWiu/RWjrvjShF
TGlaXruRGKKFQfxZuVaZVTnQ8TGiPO3+jiEgVkowLLW9f3q5EpXBZCXsx+WVrMreO05CZwVy8aKE
aTduvZ1ho1+etH0wu1w2DU09QKXQjaA55JMV2JYYAmw3rE9rH0Oms5dZNOGxUVbhM6Q8OrHhjT7G
6RGD5MQN2R2IG9LYYD4/BKP8YcYJx/FoPtw/94bM19hSrr78EekQs6m0VCrNzOA7OVhiyYOJEDBU
+IFqOsvlS6nAl2OGnXBTbkHnCfAI7cHMrc9J2j0yPhwc62LDxhCFY6UpMxqtaA2+2sGKiqIUobB1
KZo15fI4XAKkKjueq0Nmq2Yc5Z2z89Mb1wSE+q/0BD9FID2ey6KdkYNSkhAXmW1B44jzwaBM2FyG
vOEYdCoN1lnr5TrRDLWMAqLq9TuxD+FV+5z06Hec6p6UcJGkCHNquC4w5B8ibeAvd9ZpbOLawsSy
WXEMO5dchFEBmQt8k7tGe4np6k8Teige0OtcfXDouQJQt4BOS01dZg9UsmgrM/lYPC4aKQ2aSn3y
QZCp4Xq/kgv4LHDlNO5AqCCZPe5IEPI3TEbHYrHZLx/btOnnNsYT+XNjB+e4wg8IdJ2xII6u19MS
2jaDDr2ckeYWMB6e2Z+JCDafDuYZF51Uuo5Z6y4adrYrez7mZAIMGjACmy2GYvt30bPE/gIEpoLz
W592Z36Uv4eVo4nrjQeQT2JZIMaC2OcF19tkTrFk9lJfqlesEIz0ZaxdPvv1iTknEFC+Bm95DLZh
ULUboSsVJdFcaKH1TOmmgJTGA5NPwjthwbCuvvBOqrxpgnd1HtnlQNGTm39xBgYlFXL2YI02jIba
GQTWthzWpBvZ1/CGbjLkYI6qLyOoKq0+W9DvlhSufwUueIzJMRo6Dj+f0H6hT19QmlvAnmEqu9J2
wpnis6KSf/dkqp0D7bXYA4UoHaW9AVfb41GLFfIfeDH1t4XY8mYyWkcZPex7Hi3LONOV/EO5CRJB
2j0CxEcaRgQ8iBHLGw6eGD5viaUtpkIpZJs95XVlkSGoNMI/IHzyD6XeeUiBP+IowH5stD8Pelim
/bjnnPkDccFCo8GIPZ7bi+xmyAYM6K68k05eryTt+AbqIwdJa+Fk1QrG0Py1djwdleBCMbZsDx80
diqM/uBszkLvcwpHSujJU0j0lvp8yi+B1jFqU9wE1mUQNz3JQO2vlU5fknoUUjdWCN4k/jZWMU7D
GyIeOd+8ONrhLsmswIXKmkX9tTP68YXX2qcdHVXjC46LDAgDgixwJxBVwaqyL+rOimgA33ok1NK4
sITOBHDrOD1EGUsMZGLmtUoGb1W6XX/gULhLKC0TzE2hOStC3FGSBp0Mc3+Jmy8fypWrPdyzawvN
W10cQVcHpymb6VdqKyaAiGad/+56GBVJ8VRz+Kvzfox9DvIbQzI2GA19QejwlKDmqgyORXB8/1Oj
JrLB6SVqEgrrts6NkGhcCROYrSLXO7Nxf+t36idnR9goOU9n9Sb+9IjmunORj75ZP+rf1C1A98Po
43Pdn2D7mtcznMpoe0Kl1g0tHfjztARHm7QA48eeYoDX3yc192vTuNUR1O1V3kReQ6Iz80/nEu93
9P7PZvPjg4kE/eU2/td0HWmvsTEl3MNiXRpFQYWXHGSjxnQMoSMXclEBpqS0sYHyjPOS26oedGFB
FxbpSahDOPGHUR8QzX20HEkdh4oEJC4x34f7gjuhc6NfOb4X39P5fyUoOIXYreEYli1IyDGFTr5V
5R0V1rG9rYZ2WtDMbmPR8dUi0ckIGHXcVzcBJxCxogjd7tIZfAo7IaW0dJADdrSozbjh6+zq8KkT
RQd5rH8U4NzRuMIHMvE6YA0/IIQJ6qE5ZxHGgLeGFfFLyWYofhOcxSOXkKjwCryVa5WhM0mSQHI7
vSyKkBM9FtBhwL+jy8rxyDzBHIAKq5cA8gULZiP+YRx6IMkL6rqFd3pcr/M2j0KMTPY1va5/rKb0
gdnvJhwuIFelT9HavyHVs3i3ORT5qVkyZboLXjlZ1MkShiBfWXdcoFndl7+D/9P3kgL9WcSctAtT
J3FDqJSFn9eEyNCn/nh3bd3m3IxaLW+GGj9yUL4RgBm404mPGbzE2DvmLMSKRpEp7P3+G5v99zNQ
PVsq6pP+uH+nnQsNWKfOlx1W8e4bH+x3gb6vah34EUJxzeardOk6O88P8HsM4tmkM2Zm1zMmhpTT
jjlJPYcrZAjOAsQm5mqCaRqNeGkiFL/EkJgD6bsoOv964uYC+bHX7aY1D+zFHa+/9cGUhh4J67xN
WESzTDCQusEwjVEW6t9rnn/6354crMjmcVP36LnisZ+zwfsTXmY+kMY42PpjxoZRr2D4K+u17up8
9EfppOiS+Iecyb7UcKt3SKSkg81wGRIcrhsh/tLaIFPMS77/jEzzD1/VsNkSTC4rv+/B9iLNJfm/
ITv7WE59Y+VEEPjKXLGqrU9fumqTg/AxqIsnJofQ+GwwEHUjeb3nyR1cnKSx65boMxfF5MKqxq1I
+UMvrfyuXjh6240OrDJWBL3kJJu9VZyU8zINxy/VoVfDvNkT+f337FA3wE0FhE7W7R4OGJSawFYR
IH4T8ytSsmNa+DqI6sOSYYis07DXbbmrrN1D1WOfJ9o1bJt5On++FRdnm9WaRp7/kEalsaP7DgWM
ob73szsXeZ2SomzSAO0vDBPzmWecerCC+6XShKWyuwWeY1RARWX3OsXpMy2qyFlWQSV5XFGPFvbb
jlKFVUxpluUrAJHYbRdH6dnrnRj0FYo55yuEqb+dR0sv7HlK2ZoChoQzJ3xRBUw5WFsMmyplz44R
nTzq9pZQ9cOq2gg4E1WjPxQnTGxzKxY+h2cJU0WkyfmqUZ10bMtYfVwqXJS+O8thzDTJd46tgNTn
6sUz62NzSHsmtaWZczZRrPzFmKSFOl79O+TCX4fay6XoiiHDA6CVBbB7+SQWSQQwirr+lvwotJyt
mjl2EEN0J+FDcQ74JSwVEl8bAHZGk4lvR3R4PLMOlo/xZcxlp6bE3T2NwbJiDvVjnSafZMBiLA5t
S04wmAGmNlNeW2TwwfBM3w4nnj9vMvyhehkmoaO5KrVtIgsiGIZI5Sly28Jk+MmkGoH+GjKxwf7T
AOwdNt03Wq7Og9UWqRegidBXf1SnGLQog+XWkb3uxbaUv8GruEw93xQDeCFXG7nhMvizQlwsvABL
bWT1EA9p8Am+XCOnrtB8ZlYhkeLZxu1Uf7eAyH/GRpmshtWnuWgrQFiORR1noxd7WtYg1Hfs5p67
oPNYcNYPwb34XQ/j0iAzq4n5vYXkm7netn+Gb6nDaNGa8kxOeDbvnbDnXpJb5Wj6f9pc9j/VwlNo
nHaG3E6pqVvuSbhPoKh8ZusvA2vvClanM2sp18ndCHzNJm2tUX9lRi75YuPGMKvJBaokyPho4dt/
oTAF+XkDh81T8UXhGNeSdTK39Imk54WGdkWfd+lyhbkqeUyv5EDBmGIWd6vPcHprUHAYo1OErM1f
wH6MPPbsVMRvWtSMJ9wrY8UZwp51axufcnJbyVPyxUjhPEPnJu9FoKJJu74bjfUAhA1jzzZyPfoe
trFquXqznwOKTbRuxymVAS68IjVMJNhv9jHWmM/tAq3kZlNms75Bz7WLZN2HQn61r3FNb7ZFMsV/
TXdJ1X9hyGpwe8A6M416KazKLcpDdRyARui8Nl1H6qeByQ9HX/2rRF9Rwd/kCvG0eZC6ZGvzwQSC
DXuwS4YGujhjGFXcbssMOCUyGhtnji4rehd0tKlxcPaIgG7mXJ2ZXhKj+5lUHeYU9EehxDGV1Xa/
f5vv7lM57bQuhVST7K5azpiJPH952HY/Z0j6A+MFm1hOUVFwnAaj0RlDZ3MFgtBUiHBGJ0Ai4I+g
m4cGr47hM0DaexkKRTKBubYaQ+Q+4oiuxo9fb5wZ+uLqFIe0XJ63XTy4uDGjItU+p/EYXkcl1879
umVmFGedjKiy8Lxssw0Xkbq214l6cznkWNRtrb7aaRJuv/mWZuWnGv9Yu4WGVTBdpp2dKeKXStW0
gjpz95DUmG/o58qix2fepkGTc5GLO0yTii93DameK1e8LeJ9tnih4jkHRqZE0qyE2K6ze8RqSsnU
/e+Ruek2GiIY8tcuU6QP0kE3h5iRy5qf77JS1YVNsPnoKNZQIA7yNeGBCTqvoz+XXEI/xKRBqojM
Uqf4fSHC2JJ0HRRzDATTgdf63iNiOqwwVDyjVR0IochJWYH7MV6iuPR4FykVts1W5Lp0Z5iQfyif
ZUi5Dr7HQKNJqdzRNumOUfL08u2JmgMnfqW82KZ+9DFafKJlpCRvQlDY+hJYkztap1/LAoImRCwi
vWFn5lFgOs6iOMOE+1ICYZ4EirQvQD15UbBBAXA5khvDA5s20cimJqkgZ51yTYPvA15NG6NMjM0w
5MFIfSF7EVnkVFmwmVWQ4Is7lieNU7CJd9+3Qk8WdmG6oCwhRfwT2Bs0vI3FbDHADTjfh8+Qc7d3
3Oo18e9DsCPAemryFzAfFY5GOvZ4QMi+SXDmtlYyc1vQCzYJ2LyEzNM1ylNVkHO5YE3RLyivhaRc
uhM1Rz9vU8MEd1kJgRslMlvsQR2gbXgnWVTTuVl+JynsZm2rrKGCBJlZNjTL83ex+WkwMCnW++gE
watmgKSYCDBQJSL2ilBniM0x01RlC2SHHmRH7Tp75YgpGCoVIjgMSIRgqNfdnLLrBKKYdo609Lj1
LkK/CuEMidJbiJtB6wQpWl4jubg1CUD4sUvt1RkmVPbebu8fBHxk8D/3ohna4fdYi7vKjy/vtMrA
00Lwc6C9a9wLm4GZZDj+7Zxg3uNsDAiUVj6jhG1AYgF/ANfPhUsXC518kaLefb6seJlvg61Q0RUm
yA5K1iQ/pSqv9H38LoZJqf1VSxtQaStgqXn2sWL3ukwize0jjdmUHerwkclvIZ+qn9EGiHd63Kbq
dVliQeQ12OBTYf/GDeXVfRyv5NCaxVpolIo1XU/mmKtg1pzN/7t312hhHSq573/1cqpa3JhrP2of
21d60NJp8TvuGhFAdfNsDifGcaeMGPYOcDCcDDsxpPLmOpnwfT+iNY3GDQN0CUFvrZAulICZY+db
zMTzMEWXVdHzpPV+h1faVlmyHdf2QJHtV4oIU5FMH3c4fwqVJj5kHPzTEL/Ot2xdxTMh6hGPJO6D
u3kyfUIkO0NUWwCrZXLG1XnvICF3crUsDF2y7eOucdbAcuV1rrmJu/6K1VDQNehWMC4qNv9FB6Aw
ryXzNnUcHmbiUjTdlCupXfdMu3Sle/GZE1RV5hX0ExJ3xqMttRnFPvUsgFfNHC6uXNN1fe43O0dI
yn9CNqt+6ZEn8FQW4BnsPZCqVxixH6vd2ogPiCwcURuKZJbujTKAda0+loOMljqBUKU9rwD5GLZ5
Ja5HxjRFTh2/nbmebME2pC+Ckl8qdSa1nNZed1Wn1dMymtwzt8bIprkAWuaHJpjWfI/GWYyCeQ6Z
4siIG3S6oWbZRIv7c3mYFGuII+GDsOd/5neMoao4XgnozNp+Qihdch69WayKF8epi2uxzvcuYCLZ
sceCavRTCNpCSkHhn8jCvemBjcYKMgy4x7OCwVtMjxNZz871BNtx+q6cTPL1HhbAYiRA3n5Xf42H
E+Jau/K7aXU6gwjZ9Mr/xIsNpV9GXE9yPrOBlOu9EXme2YTqTweoFz7D1MmUWp5N/8F3PTye5oAP
tBpWfmv8eF0G8UAEV3iSb3vmEeDPrUg23fIVE6Zq4dsZE2c7HdXoAvpi61CnJ43lSqm90lF2uzW6
a6r4bWEJj9iT9chmooJJkJI3NDWVcP9JWB/HGATmjpv1/48Jk4lHtEuCTHhbhSc66N+9IaAq/zy+
BhKXUnO2K2oIlmlUuiXG2oDoxqEEPT4qTEUeLzTh0QEXeqfQ8Ebo/4vRJqV3Mk9hahsFGsUG4HNh
6ZzoucOcyaUF8pHNMZr8oGy338yAbPw28XC/izwgpC9bLs2S4cKw7if9fhZGDXZheE8QIuYSCJO0
50Yh03UtPG3PU85kbcVBGb0hM9hnIq6Je/bztgdXe3tjG0L40+3mZNft/c+f7zPJd75TanhlHhZD
PxGnedG22w6SsVo08IHWpsbPONNKB8KncA+23o0uY6HfNZZzjjDPz6uzlR8hmSlBoeiXe1p3gWSx
CdWaJCtFqOR2IjBoIwJuHIgmelxmQvaiLHpE6/ksaSlfteg/99eRvhgSwxKqQZ7C8uXjd1PJhVq+
4JMnVibthL732IpqEmSrLEmnsJsd/GenGuMU3MkHiVQmzyKpeFqIvHP43kRiQUyUPdauAh7knu2n
5NHiDWuVmLVxe6FZtP9db9ASDp/2rX//ubti7654kFTaK06YtwuqD1f9MefKs2H9HRAQjksp1Y1F
nnyf51sPiRsp5kCTM0z2eZjVnYpKBB9ywTB88lI4ybiX7kTIjJnYfJy1bnrxSIi4jiLLBxoVNmQE
2GG2vwv6s7iZYaDswgLw2VLoeSpYvIYlK8s8u4jt/hD/cpE7weFM3aEIVB2ZpuW+El/cyuUy1h4O
4rmNWyx7YtkGigPYR8R6b5z7SW/P2MfRbv3UI2vvy5JZV3oVpKNCqNF+UO+ImFFZB3e7ohxqia1d
q6CzXM5QwNHN5TE5fELEKfWf+PiASbcY9iHp9XPE409Vh6cnCppce2gvUsm+50rWgIrDE7yP1zG8
aOLbviQBTAEqzWzWG0pnh2vPqHKiOz9ImGZ2Txdk05msFw4aG5ClNxdo1eQkwGkPRSFUc5Mn/Ki/
vLBsWHKvmjcqrvLQzllu7cLU7Og7wOIeqY+u9nGJvvEtmDavuPqWddRpfIDD+sX+WQTHemxTyBoE
XNbyd4ueRr6VG3+3LsOUY3y4IwnspGfE8I3Ho8MhXRC5vVrZhtMTF5IdYO+3Dmtn0Gn3XWEqtIYB
8OCiR9LTCSS4sGlUAAwNytYjxEw47gvHm2vNwttPw8IY0WAZ9iSAjgXR52p6sZYb97dzfIuPz+K9
Ut/NiYvC6CmQvpJpj9uGdd03Iw87ZQgHbpWN+E3QPsrJ8im7NmpU4V8u2SrnYDcRjMpeVCd2jXh5
oD+561SQvcxFRor2fqSXYgDU9iCkANsYlQD7n+rUL5kJt/ILVrdNxWEmXdHoJjVjV0y/7ZIhKxmL
tmm3OQXVnDHtwfsThABY2Q82tUQjlQ8/yZwPlhkayFhKDpJJU7SfHToHHzlRVsxb5oYYfJ5WTQud
PBPWx7KY6c/4DHyQl7/U+1OhEyLbxYkyBbD80/bDeQwtAiinEBt+rcyYVCsSvLkwfum22lsS5lk/
4zTvLd8/fPPc8CK6jeoZC/98DJ+a0XE2aIKI//WNeCJ1F/f7xvPWQYN5Illa/HolmRkHjspf/JqA
lrgxII5VqwiI8tjuYljqem5VA4sGgTZI3oL4OtDiuEdNzXpARCe5CSNx/6ziMWf5HHrB5r+o9QCG
zOUz2Jui5lC4x3b7dTr0VAh4bwV7/Vz+R0hOuzu12E/JJMByTZRvdhvwaPxzZTlHramB4LAxQE/z
bZ3uu05iGrAQThzWfEdr6ZA9BspXRF6dAHif0Tlydr1oKRoTXzpbD/JxlOlR3jCAenh6EAptXz2M
zV1ymYWxA2dvzzpAEe/cp2OSu/enEj8kR8/PXDeqgF9bLgQuMXXBkb+wKTqyYU1bXTD3Uv/w1trp
lBT/YK0qr4P9hibTluJ1xCP+j18qxUztwjaoAOL1urL4wbBNPvgjzYaIYSBLo9SUO1Q/KM+x7SLF
QbGUtYnDSVmAANnQ2nnLEGZMK3qNBtbXO7DSzeSWBx8HRo43T8AS05WZCr88DBWmtThd9mELaAK3
2fH4JKOdJ2JMpNYvA674bbDgFqnfycjXCftEw/CXoH84CTkgseIfMVVnSJCfNNEYKpF8goqWCR+D
WCF7wvU+A8Lf1XnkS1dwEQMOQHDQDZK6SiCni1qPKbPEIlW/LrRRnOlcQRT8/9pOQPOs1EquSkJi
wRcGJwAMt/xYzXG2nUH2paCQYHLc1qpWFcE6bbtalNbealNWpf0WnZZMJhGFa2SlsjKGmHKemwYS
m5jcoVNEGifqgKaDupJ4f9MTy/HFaX549xYbo23FcgC1P2m7ZymaHTwBDf21EbBeegT3tQXqHQjd
ukJV9wb9C7tXpQR+EjsLZ4awgNwLfXJ4+Lhv/V1sW0n3wmVKLrUeIiKEJYV8hwB+Fj2SyFnnc5my
Rxu88NejjjG6JDGqtDRFpZxMwlyUS+z2cFsX7MKFPNuMtbe7K5Ev3gfNNhOtqcwmsRR45zxocZ2/
QGU54wSv6jHJol/yp+f/QfTubaUSYeAmwMqkd/fc8jmuDtkkOcm7I5xS8z0GHm+UGEnhtpfzyBvq
fqvZ4h7vh7JrzBUv/3N12JGsR5W+N6GUjbMszNZTj8cG/sO3jjKu3MRGyQ/yOwQWsihIOYWD8HHg
jMaHzrbWwptgdd0nnnxoXOLSLQZyL8Ewm3CBAua1rmMLuevcmNmYrNwJYlE6wNl7Lh/p2a2TGGS5
DWvm1Kcd/U04kNQvk1OODoFf9ZTBd5P0xFX9s+eNNUj2rYGjdoOG1fpi03EwO+Dimy7wyu7unqTc
EoGiWdF9OyGDaeuTN03TfWjcWYXMhSx84RwQR6ogEIHl+ssSH2uJJgE/rQWPLmgLYcyhzS7lxZkn
AkhK2FgBDUOaA4ctKGeaJCC8seopeR+WHciOSlRFFpfxKDodIBdp80WD8JEWKbA1YcvNqfln2gWP
FyjqGgZiDygmly+7bHbl+7gYDpGXwA1RwVxgEvLCfLs9La6hS9L92WT/p+AtGR1hSmo7yOAhoHZy
9qegGFxhOAube3vOKvtm+oOaNKTLsjTlSw87+MgI1TpCKwsplOxybG7ilqD7k+qAS1NyYYLAj6se
IuVza79qMMY0ICcoh6toseaaCJ+joaW4m4oH5+QEbecch3L5qIFb99ENdDNePjpALg18vX4aoXHc
h+YsdwoHCdpY+ta+MHoFDcy8fZi4w7PQTAMVGn56jAFdlV+h0ywEqJVaAtKNCSnGmMgTDZFHSVpm
z0QkTQCNjSwtXq0ubyCGB4+Hvjn4kgU2GPbGTTnfN0C8JZY177flqDEF4eDjompilkWAIvKhI/qe
2BxWdfFY0HKB9PcdHuY8fYsBE1rSYDILtHRTiTPovjEJ9GaoP5FnOeYVtJ8d3I+UVShXHNT1HPgS
PCWVJ22/oDNSyirJqpZ/gTpBQtDKCEIovi5B5ShSlcc5Vf3tR4EIQrrLjjdRTZFIMVC8La3CWWkB
/aM+n7yMxq8Iqo9GPXcFAzXUWRW+9aufAeTbYxFGtPYismJxw82r/7JM7uCSS9Mua22j0in+L7Kn
hwDsg5rHTI8IGeWiT2tAs0+u+t9qEVs42hFEN1qTijbTsobj78tSf/2JAr8BVUBHxoRa1GK3ysJ/
tQh9K4FlrsskxlzLOXIMZx65PG2cQktZVHJaltwRwvWIU27bymybKAtI9qTza0dZZJ0FJHiJJ3y/
zj8/zO7D91YX1JimEkzBvbS+pZenLwefSoObmXjkQHkRedktUX/6I8ALYOBsWuMV7CuJ1Q3WMwDV
7WRb/rNJg//m0Z9D9zsSNXkLtf+rJVm/6s70tNtYZ6ds/wjLfJa4G1HDznDmnqQiP+BIzzW5KnPN
P0ujEF3D8Npf2jbQ9vX7S+4iLu8QF2ayrisJVmbCNrANvmTNQaesWZG1Tdt44ttam3Q+4idBzvQ/
Ymqtgobl5RHvjZFufgMr0KkXEOyrSIcBTL8DUn+MX2g3PiNnRX6tZrzvbNdoGzp3W6kori1TT+yG
Oo1Umz7RJwRCBXjrDooJNA/xPxxajs75L0/xgGZlJy6k5rhNHXJdxR0E5m3rbcZY6YYeZGE0ujFM
2gLLENKwjnjfLScXyCEUbk0i9+cyDtKmWTrcu5MXucgisixyHJF0Njfdr3fI9KUbFJuSjq0uCXKP
tci1bnvxoF8CJ+UPD5V/hshIlUOfQU1Q/0zcezGlnp72Rx7x18OG5WssHRyXXKNMHuJO/k6QlphJ
1thGTFXKAiibI+SIo5EM21dtVFRkLLLbPgv9rcAdq4P3ccuCTJG44V4QON/THI7XGBj5p9dMPI0m
Bzz5LSRRW1N00hTkEF+0/Ks1Zvifjw9s3SmamdUp+j1dYACuNVYCM5Dd70KLnF/N31qNYxwjFXvk
O73yovq7r9AJuOFWSMiFK56Kzjm8SuH5/OeMRm47NmgUrXrkVjjv4Ij8kHPMiwNdrMvFFO+5B8Dj
RHvrSuA7G0V5HhsloiLtlpltapG1WC7qx5P2WfIFk9Vqf64DVqQry3pNfiAva1n5lM1dI3atLiiJ
DcfMJb6w9ad3EHGPgvghq6cEROq5c/zpK1/1jBV6MKjfcX7FBvQBWmvoE7GOKbF2Ete6U76+Z8yU
u0tArsDl0KtW3iU6vUAjaoH8DwSHI57GarZyb9mRdSFwWPvJA2E2zbpVXlxPktQZCi7VYK8zmEPE
NywtsnSlFRyNQLXbvCydVgbTP0dKFrB1hc/ZpPcZ5wEqDu+9UP+3nVKIGrF8aLG2A2mKSIQ0iswh
+LYfXSGrt6z6GwmTaobvRaiyBXK/9k81wMglMYqw6yJ+WFfnLtzno+xxV3/I7Af33MgFABAaulsf
1ClkWZEJsBY5dVAoJ1Z0wD46Y9Di2cK8J3FOZD7JqZDuH8KfQwvVdX8YCTFaYX6SfSZHNg6h4bm0
R4cCg4Ux6Yx9Q5B8Ybv/8dC9zpvwW9Eqn6Xs5t+5ugl3CT59knqxC+4zkSoi7psA6h1AeoPjYhDi
SSB4pfL8BGQkezNts2FJdT4O+OLbIZ0eHksyHdYh9xn/BABgA5smQQ+tiHXEBm7OEHizqZXlDXMe
e9mHrJSNYBq28Ult683tiYOk4kI/fXQ1vUF9G/2iSZT1vjfIUW98Ksq02OuZY5YEHCvKfNCd2zCF
Tw7+mJlvDZbDqn3/yFWlyikMEErAe7i/WqTiI3rxqZ5LD1r44XwANSF8TKVozaYydI6F8ZQ/t8dj
wEmH2werU9HOAuUouB9MWKffr6tfr/YorR5e9KlbwfCdlXCBypyQVmnhChIETycPQNV5QSZK949U
7QJqfc3qL+dex4N6sLy38FBV8ubTuI9H3ll4hcIoA4mqFxJrS/0ZSEFRxQ/2svGCVUBYk/HiErBo
jw50LwdQ6NYlJl0P5e7ixoC0Gk1qNQIE3M0Sko4S961dmXnFT38Unzs9ppSx1oeRJZqH2qGoo0De
RAPpYFgDkzcAXx3DSETWmeNGC7+iiasuiKiQgQZYEFaIDBMWGPg6e9vzQnj9DWKKbf/exFXtwYoi
IogiLJ+WbyQStOKpGMJjvAAHXO8E9G3au09gWGVoAqi2IhmYyMr3/Bp5OPYJo49lDK0w38bJaA5N
Ou0cpk27ijAENH8otXKaGHRNo7MI8IkNbX1VkyDh4Nagw96csFuklJJqXWDxkKXCFKymcu+MLzFL
SjGdaFFukwKiWh9xpnru1l0jpVq2qFWc+BfXvb1+W2ijMghbqj3CF+6IhV9Feck8YGeyDNTnemx6
9sfOKvt+bOVNeK1i7BDlpUKFgNV2zikVnsyfFP2IyWnBV4SnxZHrnLfx55+Foe7AkKNxToRQvVUz
C8OndxU2RK93UbU1nO3dsptT5jVJdoWrKseIN4m5K1dfbqmzeIsddddGv9gMxC74vjU2l0TZuHHd
RBpB1MLdDwvrhrdkLPKbMtRxqQ/PTUy1Ld7nChumub7aWhXEXGycIPElgDWe4xIq5tk/Iq5RYbkC
i9YW4p4l8RH2wLmA9xRViIw94QWYXCmknDtUbq+kgxPqj7iTurEegOwYmqNT9WmaRes0PvC8wOae
8z/Pqe9XyikCJKFKW8By40hLw9Lw3+JpDoxx6wAutdXwii+tgAaVJRvqDStcyCEI/31iBbfYa7Gx
84XCC6HCzhY62dn5KLt4f1FY4Af8uJCKPRjAfvV0huxH0TZI8amhrhr3tzy5IH7T04Sq/XwfZGW7
aInmLa3UC6stPnfYm5RRq9KoMDWv/eGrLnEl+ZyWEKwCQfrE60SwUZX7QvCBQg1nqzHss6frOkSR
0IehtHyg4FBvlKc3ATj9BQKzhaXoECSWpY6AjY2QhkZ7lDsnzQUhDFdfhr7yRC2ywJquZaexbGm4
k3OcfbGwrhNUTSixYMHzzh1Cgo0ecliI80w80bDybW1Fc/oQXnFlG6noRqOSf53c00fIzvwicBKi
NtueTrzAEuJdtiz/7WYreoPsT65V5GCTvw9xD9eqenwZrJSHBvCs2KTDf09o9H21KwA1GKszgRZY
cS06FgP9QpIFmWTnSWsYhmsRqUHqBnvYv1AicTzm3+2YbVPHfkJjxeP3e4OMzVEJBmxPDpnqeNRQ
ew/Dh/5cXwLz+XBPJ5Thrj4uwRp+ljKf1dvihN5/XmaBZFoy3JYIYKHLhr99hMPPsdv/0ScS6ZIh
AhfH4vHISkLP7wf2agCuWimRrYF74mdlviwc5n+zvi5LK5NpGoX/mHE2YEhy8ecr+q+iRQzDwUmi
9v0j96kCMbOIW58K1koi8L/MVw4KwJmr/OtmDJ9Lle3tbulHawSCQHxX+qlhIknTHXPv6j6tDjMs
WNBS77ujh6nTrfXk2+xhVvXhNK+3CQHUoVj+unTMeXmU6QCJkTYaMfFlM74Hs4Xitfx0tBqEGx1t
O1WJqlvUbOsxwNjKmuFxAw6YEGzV7J6iuhOTHB24fCt5LZ830+gPxxMZGsbMegC7TSKkxbQCwhTu
XMH8q3FmHExS8ZLXmQWhdjfbNcQJnQiuZeHKQutUWdT5eqPSw3VPDodAV3hDVKIZ6m923r30Gnee
pEVyJOm/AVWAN2AgB1SwcMC3rXXEksgErxhR46P8KyoSZMHqfTVB2jnfZQTk5R/l5x7NmarB4cjc
c3Ucho5m4qyBtxTn3lVB/a7HQz2XkoYrzUZU6g9FRMpLkuhAeFenJjtAp4MM3Cjq0kC73gAsWvne
qIQo2KsuFkUyorIZeC1J7XjmrZQI/v4fUp0xYeO5ASBlZXRVW79SKVg3e0yvEoSIi8Q8fBn2GKMz
5qtq4CFAd4JUCjNd+EnrQ6flrrqw63HuKFoCVXCdXdmv0K2nVahQTFHf+W6yAwdzJcnXO+1T3tQ8
NUx8VG/idhCybpZYuc1Pu2ZmG7QwFtQn4D9MUEGsn7oybwx8C1narQ4s4bBp1+7/R6VRF60X97Gt
FJ5oBzZI70u1JNKmjmJiGfAZiT61caT83aF2lKzwjRh9qhm8ynU6sWWQPiS3IqGsks9wpOWfDcHL
G9w+BMU/Z/J70X+Ij7KB11FjqSnGZaQcs+16E6b2Etvujsg3EX9QXn5DPocD1WdmNqLP33h4O8OJ
EniH3poDarOFHNZ9NTw96pMCwjfwOHsHqe2oGLyNbvnwmKOn2d8E50yCDtdIB15x+Ls2KRJVj9Xp
cPSBeB1CHgZnPU02zWAkmC6dMR5QU7GnJdtaQVVnbjhUsDh8CF8b6iKdsNIsmO2tNATv8oLszjBM
7LiNbtrSfC3vG3HpK0K37r1CICnVZB//6EtkjEk/9A955ltIeEz2FfWHuWP6M5W8s5DnByzkMFhh
TiSKgdFX5Ms4mowNyhJ6nJenuFgxztQDY5lcRPVGNMv1BIv1HyleFhAmJWIKpryPMMN5OEqGtGYb
AE7O6DlpdXxHKDQvHlW83knDQIFJsnIq9QsxdYEt/W5gWXZZGOsG2x06bm+vTsDWS+Sqst6ZiTAi
+MIedv+AMoAmYsa9zHZ94yzry9vKp/jbUa0hiB8UySClpfFlqPXaQpu5VelqNblA49ankahIvas4
PwuE45Kb4/KVg56G1xjGtDsprJN5PDP8BXly99oyauNyvQ9N3QDQFaVAPiVP3q8Ha1jc/41zGyz0
F5AFiOC5rfH0zNW3Oxra6Ov7Zb1FbndEI7w76UXYUjYsMaOSKsCa4rDGhaiamm1uyU/Y/maMpzhW
/67n4rw0NUZMnlF9t6hTsyAhBu/QR0n07nuQTMXetEZxbxJVz2gRmUrKfpsdlxHmgzLBKRlmMQzz
I/S3+njJzvqgrVIejrY8XIauDb2ybNOhEZDDeTPyrAFmCAqy1JLBuGkDslajmyl93oiJQlaXSLKI
Ne6kTAt1TmgtsJgVyRwc+1lG7UjWKzLMXKqLmwCao4X39BziyhlCymLtxajrnR5LHlPBMIEsy809
kgzwsjqInO/LPxdBbpsW3ad03CV68IUl9aw5lf6M//MTll8hEHEwhJAdGzi4Ir+tCGQee0ZcvQ00
nlSdRB2b76D/eKfm7fFjYHgK5PQQsRKCvDisGA467qRg4TtmGiI767hjBMJUEVrmiJAdJTZtrLtv
vWqv+0ANVI4UX617M/hnsMV3yVQcZi6eMWS/37WfDo3AwQJoHqTnnRZ60nA25DtjmN+C0t+bxbeY
hAMZmROIAa3FHE6BD/pZvr9fNI9a3aZ0jTbJm4MSLFrH4NPn4KXr/BSDhLnHTgBt3Zt+aZFZot9i
jdk61OUmSqVPq0+xKKjyJCsLSxhbsbsQl1yaXE9sdqiRObex6MismxBEAo3EjorT4zrHihhLcuBh
loWuYU9X/2a0RlJjPuX0J3yW41kya0f36UxOUm12/3gTfoppveibv48kLpjKSFk0OpyZAMBYueYG
0RWbmr9Gek5nlSt9AwIl8AA43z6V1EbIEN5btBOQKxETfm60Dem48g0c1qBABoTzNRcoyyFpRiOZ
z+EMDm1hadfAxNaOeIci2opoh0BxqkJkZc5JRnh8KZ9O9kv+f8gU96xXmqw+NstkUS6/huCIVgit
18DEIErSN55hMvARv7/VVYbmQKLsOkD9c8O3lp2iWds2rcgpNM0G62ihu/PKjIzM3tVJRuOIEvA+
8y5iMLTTYKb7jGNX7HVSXLFfquWMZhMoP40FKLuEXKoilU2Po2eYxVKvP8fV84vzQPBYpyxa2e/O
/UTXW5eLufdZJ1BZKoL3v9/brxldEEcbdk7uHdXYZghIgK+Y3MDMOvqyVgtmo5Yu/TJ2aUIo7S0u
XiSypJed5xTizVNzbsCdBz8h4LYguEGllVq3vbLwlJkYezTJJVT4L7LqtLXK4GU1vgT37A1bIB9O
rwDuee2/VHAA+oli9Ui7rGd8yDuFclV1+clbIm64e1w+k8d4er/FlTBThAO49WBkGZEDhmXcdD/N
08NTZl1v2lr8uLc7dBXyqM9iFOFfcL82oqGs9WEU8JiEtAr9xqqiZvjvPeGWVX32h6HyOcQqZo4c
+4BudtcH6Obw9NsepDkPFX9yvO1/XMF38B9pFqwv5/ccdWkKKIfWPikeB5EpUBQp74jYImOLEh2c
+lQm1am2AfOkrsvhSobTLDCKN4GccHWaoqJRIPVceDAfua3B3n4FgYWfa45jWSYHV/BqW+bDsvzx
bbnb6LOedmMIlJbvT5+LMtvO6MA29PYbW4qpS7Z+WuLhYVfLNwQOCDp7+wl7M4D97veLW4SwZQZe
uTu/SdceTmK5jIFDuuYbDlejKnQtyYIf4U30kuseUn5eBCHw63roTyrvRJTz7zVNF8kyWELTDM85
8SKUk2651bskjGW/wAUxxNlcv3rA6/Yn/Z5s3vf3Atace7aIvBT2WFx0bo56SV3th4QLmdltUQmc
5FV8db+gUPfgoIdkhLb9cj5X/V1fn4XoexxTukIyK7Up5NKhjX3kJ9O9PyxRHK0r4MQ/9HhG3IX9
bJBdG+RCSmNqYB/QFVNn5VaYEgXe1D1iyFpbZD1ZDOfiyzSbbd3WT0eqeblfPGC8r8fuHtnQxTPO
1PbWE2b31i64Soq80vfTMKVToMUvBWumQrJG/yanKpnVqpVupoXwpme+rNr+0KBat1TiHZeD/+zV
YibkGoTEfjfwkSvd6gcajk1vLBkTsg/IBPBFOIeOKExGhICLY0u/vNs+ovEJaWiEQMsvNlLvU06c
6beafZWoFAZPiKQIguetLQmWqyOYrjULWa0f6e2u682mzbiqR87ZDxkg2BSVFfh7+AUOznotsewR
eSfLD5JdXl8JZLKpPL2QHBu/3UJII9PUd6aJcpN5VISwSQfBEfOOhctA6SCrGGWPiOLtb0ABEQC1
cHBZO2JJ2XoEvPzc2b2uNBwfsXbZ/A8WY4rDQL32QUoKdDdpHLUJRpAvdwwqcK3fkepjOCLs27YJ
sy7+f4w7FF261XF6FgFsVCeeG0x05oGJb8td01+uO8cNQUYozPuraAzpTWk7OeL5WrhobP2h3BEi
UsfEqDJ9qQt160oxZtOQabeiiTg6B28Rigm6zTzxGCFXj4hOG+yvDZxZw/Ax4fEZGzgsftGyFsBs
BiFMQ8it+f7yrVvlew+rcNUZCiOl9FZkdepTvm8CDxSmQu1TTReiURmEEp0ebDGWU1XBn91J5dif
spN6jLwmDwFZBX/sqbfiq+gQlpFOD23ybTlggNqvW/wzEvyNiO70DH7nuOs2Ga8Y4mQzDdIi78Uf
MsshkR+/jIePMucRsM7H2yKoKhBJlduB8Eaf1PNYo5ZdRiUOkIu7UpmbJJ6UzajvArMp9KSfYVb1
mDA826ljcTSZlISfJt5PVaD4WPzIVJVCb+a8sexvgXmgvC/+Ko101CGR+xskfBhIvOzJ0Z/vAGqh
mCzRKmQzMxfJCOAgIMsy7KFuH1HwFID0fFPBv13X9l2tlwgSpzYObvyjeedF3FCtsARLyYFw/fY0
8pByAT0y/9kEP7JRjySm4V5341CQA7RWWuk04qH5AwGafZ0bCbp4kLRI28FFRMe1xlqg1VMFueDp
vIvAj8E2urYOz98hg19+VFGUZvneW41WTNwzXJcUbVSHtYhhSZsZzT1y56rw4H8qCpahtqSZDjjl
RAxr0+mxXpiQKl3G31PULC9ZwaBVdfctO8Q3NKJFz1qAgQ2BQtuv4Ng1532pRcZmbdVLpX5BNYth
PeULQLSJgA/auwsbMlfPEtqzdhCvznFYGmAtX4RRDT6o9Uvw3rXAsmQuc30MK47eNh7Vm66bk8Q3
jhZYIo1XKW35IuyJPpnd1ApPa/pVlJVxhl0w1Qi6drjWNX/XZSa2vpoiDOJ84YTClUhFp2cRya2u
NdhEIuOfr+Jssv+XbpH6JEfjYTfIODSDyeg+aEPmIVov3JuhHo+Ij5sjxqkqlwYLA98x9t2ebJt9
Bp4yDlC8ktJ7t5nL8TXorJhCpAktCfWXOBloDLMuD9aLw/hLPSgWprecBjcOf6Mr/Bfny6BFrHMp
6lHsmSHud/1NWoDMzvhBMCeIUn3wwsPoYsOhUfXhEXs4CifITmATcCZFiBaKVSN9udJIhzp8ISes
tBdFP2Jed2j4ZKeqswOd8jUbKCldArSuWPx9R20WaTFvaXwzDWw4s9wDl1+D64q9jVkjsnRd2epF
Q+bbU3vhvZ7U84j0X/+3rvjMDTgeaCRjJod3N/uQlC3maJD+Dq1eJ91/WRcBN1XdKMYoJ1fdsi7J
fhjKqvqn/xDr69TO8p0RfGWnP5uBeAN7RCWcH1YJyWWNqB7ArPRvjzxp2Lyn0HgE7ljq65h93DdQ
gr5T8y9Ms1+Y/3jQ7hJc2upa8Q414pZcygxCjLqcBf9XpntHXXwQcoljbvl9sBXkfxM2ZVnFkVez
2oaXGlfD/oBH857HLB19LwBzKn2IvIkZEaUfWV/Ig75qCcndklW8pduhvaX46e2uzBI4X8UZwD36
JSpNfq973dBSJwWRxj5VLUpOj+P2GDKCfupsYZZSL5UUFekEdQe71Dt3WX8XrW17UYLyy388pqJT
+AGnA6lrpIH+h2p2+YV7SzUMKqwVQEVn15SpqwOurOhYsRh1mHHAubBcF1H5nczJKMHyJl/hEH5f
HnPP9pRgPN6XZKAYs1NzDeWL6F7lpecc5GCK3ZVQq9bDiKkRlpP3Kxqd8r6ZcTpJzFo2vWiWMj38
kRq7t7fX3GS8Qx9+HBOp7VLSFYT0AOhYmCIXWvIHMWN3f0j20Lle+poclt3IXdYV0vFlM9QP05ap
Z5tVl/YTSZ/rdm3f4R5PyR0ptpQSaZbiQZr2OPtqI+XpwNQ3Csckfzg8N+D16W+KaJXcA/9SI/ig
KtT5NTV/yFWgIhJhEtFYsLTkwnQHn3EsgVcytCZtAKdt5pAmo7c7oRQuNLN2FHe/esQeTC0sQq0d
I+/zGdSdQCjYPTdeYBWNdNov0zaKG4fNEDsYCGtQXmAcjWaj4WimZhuKrY9vpOaGX5Fko4XGB8UA
sfacA1l/DFtWYYjDho1XPBovGBSqIVw0ADxzraO+XPZ70h1D6hhDAR+Kl4a966t4ZHU1XQqjuPwu
/P4NV5ySvAN4I9pmTt6X22rswrKrtW107/xko2icSYpdnbFxJG3Cz8LaZOyNtf1nztzGTiVZtch9
8mnirmp64I8VmxcFMwjOykIfjC4zcTDWgjWQTzzHMloHHeRx/TruCUsH0f1VEKDGdhUPoFwaKwjt
gQ0DusRqbg3Sy5bjF4/xL2L9LuyvAjzCAe9oqgFJh8jvRlpZV1jsEzXpKDT+QUgzsaVFuGF8VgN3
GRw36xs5Pc0qz4b1Oz0hNsm8QKBtwgJ2OgOoG/e++EGlvmd8NKoK+aMNHYe2dZMTXolMjIWw9DIC
8iHIifX7sqT9nDyX0bLYXb37iROK7oKSbsdAK14dbTnSO+SzP4dikimPGSG8F1aWPw7QCRFaHYRx
B/6wetA6tvbmxcrx40T+T8RKX3qvHBaZGg9gpqLU3roGuvMBoJCidSTlmusnvxbC+ycImDpY1CnR
Kv3EzI6OjEwK9mKftuI3aKgQAPi329HqkpdNDfUYZYZbtqLWaPnuSrKhBgvbHa+qnb2NFuAiE2bM
U8WyrAj0slhVNMuc1n+Vu9xxrA3SwYUceVL+gcQEiZktTgVK83SRUA+pGB4fiwg7QJ+h9zeumP6X
dK0J4gdQvynJW1n9LSB+ix+9tMBhAx/sAiOBM8D3jqHAvyIUiFRe1TvKv6Ro/0r7IFJLHb17Hsk5
n/gEVh/rfO+LLFAXUxzh3v90TWKy+9/hztl14KTRTAGGQsqZ1E4rO8huO2Wy09jq3iMcLxljBhuE
pMYN2Q38sbJyn0ZXH+wkT+gGix+csnAeyjuA6oyF0D+/wsvDGsyQH6TFnxKBk+lfwQ35lu3LCjT/
qp0UW408Hh4KpfpU2OZVCxS0yC9ZBSCKQ3tx6n6qki+uCqn7abEHt4Nf73VDypJFxjKrp6K/2NpL
JiiIaY0rOEIQat7Ks9yLnaCLUCtIt3YIKG5+PdTR4rNAtS3MbPZik59aY0+cd3V0XPj886o3tMFV
lLPamZ4gSRU+PQz1W8wmu5z9dNU2w+W/ir6VLcAHM/U9YT2qi91+nc4p6Zzbgyb0MTIroTSEZjFA
q/JSQdO9TRW9TClaZq8t00eXKsk1PkImpgw0Yl+EpgWcZfcVizjJE58xZdy7BjEWwTPPx7eDouhJ
sFwEfjZtvuf277KdU00IMXicVTRTcYmFPfMsfJ2yeOIsWO1rXndjThH5gwUjlh5sUSC6CZ/smsss
TG3xtEcD5B43RMvsRCb1MjQGiFASzMzdb4A2gbYd0RAwRE18k+yvtmxgu2OMb117yqTsv7x7pLLm
eZdpQ/Yut8Vt2y+KEPRKWSXw+TTRiVW88buSIki4JZLPRwf5UUNENbqmGfNV4OT/cnzoo9qXluGE
6rmcdT8p0DSMTLlOjfflkICe4d1XD1xzWANYeljS2HzGQdxQ47dP75dEiU2mi3dcZGLxxOSRnyBG
0zjrv9GqXzIAyQYqp7UdywFmbe5eUkHlQ5qb5z/teM2ywpnIBnCbcf60PBdorRLr2wo5rNS2GiG3
jf7iHYLew/v30HhVGNBgy/FfccVWljU1UWBNj87osYpE9bvRAPYvPQ4T4qCHB6blwAI4IuTyGJGv
uuHm/9bA5Zpj3Kjsw1VA8h+qcwKxm0EXcMZ+egxwpujpXUusp0eOryEkVegg3USGjsIUmbfx4Z8T
WqnOqh926TExuy7zdip1ssVdzJS3tI/AOGK1MDN03j/xwMTyqTZkkcCd/elvg8B+ho9aupHe0ZQC
I2jnSdBnYjMkqtdT0jh3ACWDO9S+MSoOWkzK1yihOHQdaYCCr9dfKzTLAH9Z1nu5kRr6qNGbvnP3
TtvbGtEhNnP+oeWTe9gVirJyWdAV5EqheCTpABXhEf6MU0s4JkLQG9+NoJs2HvW18J/cAsh7QRxo
YQezDd7C7E3G8kt4V2B2XQr6Ipi/P82uuC/izeLwaZCCEWBENzpygkqZDQeDYtvmd2GYK5hSd+S0
klVjPJajX30bH2EDKJgSWQUFXqDBGX23CLzzR+sUN5WzBiK5BKK9KogJtKuh6IKDvlJTMj9po5p3
rkrPeskaS4tzTvITRjZ8QbN5KecGKLgI0LHZ185Cujh3HD32us4PMQ1U/XBhwkgjHZBA58wjjlYR
yjfMWlBTNMC7APILGzWELcbwSxVbZIyKgqP9CJACAOrKOSCSL0hURb3tX2PGcCSHhAf6RaC1R8Ez
OiIF9SEbHsEUJgu+mic0HLiR8359TJ7a3lPTKz1OF3TGx/JV1chCY0SIbEab2ntftU9x7TS2o5nQ
KF6S3wZ6OlxPRC4O/ilwuaxcEG57XF6+dJy7aQrSSx8Wc7FM6wVYMuY+eoLXwkUpQrZ4QqKKf7SJ
AzW+sUMHXTFaVSV86Xq3VhtfR19KAV+Mx5EZhqXtgWq4JSWEuuPTe1cid0T3MioqFKhipLAVX2V5
L8HURU3au75JdYRR8lM0Thwe2PvKGrt4v1YwQJtBEBin/wcUxPuFzM/fg3BB/71QERhftYuPGJvb
6V3uH8oX9G8G7zrTTYoHW3ewylFqVdwlzIT7lDSgicwG8B+82d5cHWrAnS9MPNmSnbzvCLdbvEB1
8lY2SuGS2QskPjv5AcvuBvqS9P2IiBRDY1Oa47/HOkFvlPFUIF0MS4LS/UhF0PeuQ9c7XZTr3pQV
50gNjmOdxzxGjG3D7TNaJ5hpyjOCBRW43bqAdJjWoaUnbL0wPnNK75dUA5t/d5iQF8MFFzYi8A5F
InYOzQ4OvKdKVdZu4zo92AzLuEH12OO5MNGtYsRucykRZlf4Kgsw10g/ECfjDm7O46jP4qfVdT1E
BJtr2HIhVi2I9lPv9dMO1mf/U3IUi8fZU7fVPQtvMmOjkWHgUCj4K5ZeKvTGD3g+wfHJpDO3Vxj7
hbXwZ0woI04Tp+KrrVtOqzKzlIho94BQMSFe+8wkuH4I3KNzTPydzYHHCj10CYixUclv+7yeC1XP
30bYpAsoB2VfnSYck5/F/We1RWwP+hBqM9NAqk7cI9genbjgQptLPfUW1ROJLk2wUYbTIzEyqjaE
jQCuQN0wjRDKqpY6hl3D9gx7HCMddKlMOugbebp9qOhXFrgY8myF0R+BqbzzdaVxaI9BdXO5E5jn
Gjwsr0wSr3an+yEGUHfhTEqdo3fO6sZVtIcJwm+cWsDVT3HtIy1VrXyWTYQVSBuW5eZ9/MPRZ4Wu
Gxqo4bNT46hkC4dbjPkaURij62oNxg8szqPGqbZSdPgwvn4NDQuZEKRi4WzosS7sf5Pz36IkT+50
G/gWWzo8Lbl/fmUvq26gE2QEOmgs7zZgmiNKkAPkXsvSZRcEpy8aSn8N32rZ2fQPwFDAz6mhdHkD
e0oxa94ZQNQlIc+5dcj21jJJjR2tml2YVssLwDvnozg/sIWwyqjMd6aihex2GR1pkUImvUoZUiFG
srD8av4aPP286KXX7S/68BZNVH9ZgqrwySzVzn5RIHCkX03uo2HneIbIM4ocP74fjXXi1gDdjITH
oiRNpNsTIOcwhrYTJRRr2KdSwUbh5XLV2AQUEB2g/2az8G+9JgmGE8pzGXbIaZnGZgJITQaEcWCF
EFvQRiGBOxLyH029EN+1UFBPxEJmrGbp+ZwEGLv4nZ0Nz0UGh5jMGH/RXuZxrpjxS5lvS7MY9SH1
WT0QWooGyjqiFH6q6Q/oqGKyZ4Pm7egD/cLwczXQmGtxpfjQTjo+41XjUvMZcOqlIfe4uPHYLK2I
ZGLRm0jQ4uHo34wngrmchjWFCSvNaZutqDgO/VqhsYbv7WDShW+MRJCxodPLrTJS9GE8udqKgvpi
5ggoLa2NMalmcRLAyde8dWBfa8KNVebnSVn5oi8K7htBnLRlD1DEH9Qf8flnqBsph46OxeEeYjqv
eX7MRIkG30DvSCebc/ijdsxfOOqh+SottPPXKVMv/ri5vBOaQmPQvbtXf4IXwE9/kZBF4c1Gvbo7
A/r6s0OpQySBvxFxLd6IbzOpMdC1zVABBRJRA3GIvwfMQeqx+NZ3FdOcKuPObQS30h/vCni34r2N
RoIIMx2xyzJrJ+wtFRgeUKGVECWCiijuYIVSBa90DRWz6PK8ZIj3/ScUFg6QBF6j4ihOrraToA+G
S353QR/4AAorH1w/mG5Xx7eDsChxCw/w5FfdqgEgquOEfw9bPuUKLmRMVg7PkQ7WdpbtmSXEjgsu
lBHvogDfp4NaiDVhAN3u1sVuEua91dP6G1GZZefgMpnMldUtGroHzF+QtzoptpSxgC/sIatUQHDX
CAiDeN5NkcU6Zi0GNvyEz+1Tctw1T/PRi4JgSCln6K6tX7hTpl94+vKpLlGnQRIoIzAIRmENvAGK
1qe/QlRugs+Jx/r6ta7VNPPbdYSUAzLgzFH2WgMXbqSim7GcN3m/GFUCyur7Zx1Z7fOhn/+jfrv5
IjhN/UXbJkqlXBKAKQpH9PHLwiCH2yjAAju7t5Yx8JRBFVcyViE57fXOBOzQWUDf6neK192/GOZU
U7gSU2BSRGqmF5BpEKq67gi9MAQ6gjiX5ZE9gG5VsqRqMT3OMUwD8QGAvma+tUBp21y2u/Cjwi3Y
E6/uvg95edUZljlKDRomDe+IiDYMQOFhbuyZGMcvtZZdVwgOiTP9tngVJkc26IQokeLzC2hPR294
Pm1gpU/yibD0IoGKxZSvLRCOiTlp9l4tCjod25Bp6QtbKSjSpp5lOHrE2AdYy7YWhoMWWhEqpf5m
fRCZxTtLqRi85CjWR9g+tCwFf90Dj6yWBLIux7khi0YrLMqpfepVN0CBnjLjvOH76nu1PxFtSuW4
3XDiI3ufPfT9fSbM5s+K9Bm5lS6xI3wkGLjoPlryuqi11CcqDkcOR9CEz/I3/2T7dalRaJ4X6yMC
zRRcGoB/O5/nNfxrP1X1F7BKpD9mHBowBvqnRyqsD6ONvRQjiXE0LmzrAPB4Hw1dQJIgqL1prUK5
8UpEUdrlGyvb7BIb9piXLCKCdIR9vGGu2PJZAb8DnMtwNvB68gXP9iORkQQbR2/QBVCMK5o3w/CY
08KD6/xfdLrvxhXv6kBVZX1oKt+CRnJgtZldXPdHLvG6ze6e+cVWBnQjs2A0oo5KwllVloNXYf0M
DtvFszSoHm1xrLhrQhHfYzf2ifyonEwkwvbgFIofcl4X+knj+yD2RVuC0qz5zVpP6zvz/hU5mQGz
hydxLSVctv8IyaeA4b/CXfMJsLy2djHVjeixKlXWD67BHoDkJ1crpDXhgdxabaU+xe/C9RDb2v2F
s1NG4S4KSmaTdqTb0rhaNzTTxvVg3mgbKzme2NfIsmICljR++6gw6ZwdwoZdMyMewAoI2P+KXVDF
AeugErk2yWVaSoothgavkXiueNZF/afWowKuUqc0sRHBtA4cDhb71QvzRZ/3jvO8VX5e+2bhYFl9
T7HPYcT54TdJ/2j4T0vGZBy9QjaGgP2ZsXCdCWZozkMHe4hYXiJcTeNJ1g3mYGV6Re/10AiPymeH
pupczl95nv176UG8NIXAmdjwkVt8Irih+ObaDvQIHH/4d267AStTregEYn+rj2K/7+ZUuQx70rJe
xKz33LmfzinYRdIDcbIb6k0lLmZ/XDRpeK8Fw3JXglaEcRoMTOAtf6n2KyE2sI7XwAl3imToH49A
S7dkwIjxN2R5RTx9l4WaZ2Omlxv8u9CiyTan7+JEBcRe5zOSEzdweTVnsMCiAaxqY0fN/to/QV9u
wwF811boqqVilxRoZEgOmbJGSNC78KQHIJUpQMabckoVXJjcavZ/rtcaMkNWcs+PbAGPxFHiSAMA
Ut2id8pQK91sqjMTFq3fZSpN0nmCsihHrpI7X/YyRCCG/hqD6w5B+xqhOYsaZSaEtlKKcZ19kqpo
rk9BV1q+6piilrO+qhl8nm3o9rs21862xshOcYXzmMgO6Um/UhQk8Rq/wauAYH9QRyaMZUS5FRs1
ccLBh+YvKWJoXK3YgkXYQ8fUX/JdIvod6qItKZGFTsfZ5toGZUgjHgBQoxK3UOhyA9GSmWDoGhb8
EC0AJ9HzutdJ5qVTtF7O61XNhX1TWjEQvuOnsW3Im79yMmh1VEyD+G/uQtme6rsgIxIZGua7sOpJ
6xePZO3v2NHjqG5P8qaGQPs/h2GmvAtcsIaNh5pAsH2f79vh1xHMbLRxoaKflMcbWbmWQo9jVI2t
rnO32jwVCanUKbOiuR5XeAIKd2hbakBsGlTaz3knGMJ1zxN7GvipTr2UnHtz1G284jUX7TlGjT6X
d/EdwHzcKM0KUX8nyoWM7RddLZm5Re30v8LhOW9w4jMXvry5AZ7yIQh+PvSHV7zRZh157+22a7YV
1M7BrEz8v543qQ85zM7zzBtEmgop9GKuhg611FHOwpftd2FOR+aSwT7lCunwvUTcrI9QaN0wAf1i
LHYnq04M5h+hk+3aaYEwHPqQjIsKL2Vs/+VIIcsxtDN2z39b90XT2DGhghPkYyzyIKpo4f5LOw6T
uAORll9fRta8BmT7QHKF8Y+kSv7TD1H7wCH4zWVt6BRKhCstUNwLOoaerK00iFk//ef1pMobnAss
xpCleyzDwrwGGxYfyejBMrpp4E8XEwFPS2OpUUS5HA15cyu/BCQOXbwD8LA9EzkDN51iIaDQ8xLA
XhFUPhE1x7EAJzwvzkVAp/FNndeRAd9GU2VKmaUsf8uoC0vtC5kGdV2N8eJXT5SmRyuEp64g5Dfk
rQMry/1svRTDrdkaBggKtAmTREcCYDw1Ko5fHum7Zv/wzQ/6Df6EhXLSs06rm5Vo1sndllwsGnwk
F1wM3UmHiLjIDG4u15Dgyf5L+ln0tqYOsqz7l03ulF2z6WSAfSw+4JDnhRzEvNBjQnmE18ZEhnW2
bVc09G/etYH2MoaclEeeFHOe7n3ZBCgGysB3PVHD5Dblkqnm5Kk/0ST5hl3b08LLKVtHlUwlCyAY
iG7PVA9JhxyS46QkZEG0zp8ZaMRua8QocAaRKjE0iDsnM/UGnnDjEy7kXSJM/8ef6CrODuDnrwmd
D8ZoLyl2gTguyKkAbw7o8K4FAF3wXEFJZug8ZfY8J9x4QddEn1rkI4ztI1Vbb66gvA8m98pTkEhP
4yCtnlXxK3rFGi2bqh6MhMrbLsNJ0hy8UoDhGY4pHiaNNJqg4a5E87GM86GMAR4OpCiES9jmZ/ea
sfx/nud1iFiLhFzuE8o9kNQfGbV4O52vonGCS6yVXn0TOFZjSsx3MBXTrFkghsCGmN5UC8/TlmdB
1ydLiqsBtfAV4Yzp26YEDAqSRGgqD/ruCYT7A6N/SWgxcYFjLIkGVHruoE7L2gOnyaQFOlhlSSPs
vZn3dtc7pnQqbsUjgyEwxmGPEiFlcHaYTRQmesB5PADCwNK17GEVHJy86m2a64BtaVRtLP+Piw4Z
1XtugbLeKXi2kpfFx01663EUabUx+xw+XA1NBdBoAmclMOpRuIjV9AG6ePoZgjrdpKoUupYW+v2e
ZefO/AIeGk1mNq8iKlEot7fYF+2tO/DBbAkqOQBmkNWW3uj/tqTeZiR2jDVKe8suqVph5w6Ut2WI
6K883CpucMe0CVSbwFDhUci+vOnxPBMPG+s1eSWv9EJ1VdxFB7JBQEQ0BPHsWckhPNmLMPCgf2vx
mWrdYx7YE2B9sNVugGNqXD2moqawkNhhujLw74daAFsFnesyVm9mpTCLTpnXcB7x7aCVPbY4gJv0
ZbvUTM1cHs1tw6hEfHuL4vSvzLgQAuiT5bk2tdStw6k7BjEvClbTQ8npNum4dZf9GudaKBV7gpYw
gPMINnYrIPctvLzWrhDhcjev/9VWkqCKzPABneVfzgavlQ2KmnXWXO0Ac6hA5gGjMde/wFKO0fPj
vL1ipLLfHilLWfgDLel+RG03SxdBGm2FpQDCbpCoEMl1dJHgrN5E/rYE3u0zDZZBeJwzOEhYv+3k
lVag+PpvyAKJQr8zamdj0eO2fW8EPRY3WLO4PYOMIVb3aKUcl6KwLiSQSgM06ba/Yh9PR4HMiDqB
mTMxxKDUevXCvQN2UGRpCaHkb3XVhxwY4VpAeJLXxsBFht0hbZrChOUceJv56Ia6yViKFpV3w/a4
V1R570lnj4GfOIoHfAhcJYs3QcnyQGhthsDzW/TVaLxnisfoqjfM2cA05DieH6cQGh3Ck6OvQdX+
EPeH7petZMamkey78pXed4FUMzyWd3dKsWwO5qyQKzz46OLeDQe+oII1IUtbzVs0iXIJhsuipyee
HEW3l1ieyx7DI6R7cATS/fw7qFC9JudPQS8c9WC/Ng1TDGkgKed6RvACeEX6e4FWzug99FMh00Ai
69Yobfugqb1iL3ssptGpWzgpzRElB4gcOaF+dROd4e68BHZ4T38i3PyhV58YW1EiQBWmYfE3Dfun
yIq5Ium+EI6iQ7VCEPVdhr3Ds6Ag3u86Ohq5b+wILuybSXUXeOLarZOrgiEURCZrrV0kpzgpzPg6
GNZa6sTL5UZgf5Gi4Ntt0Dg1ALqHdaqgNoZPdlSuqI6bJ+aO/SxW8ywhqms9F33Wd2beKU2dUDIO
SqOMAbjtsPUcM/CHmNQHGe3ztPmjRevoryqaTmPZ3aot9VKb3Ln4pyOnF7WYodF5DOOhBvY1LsM8
CbiDJmG2tpcZgcW4oAPEz6RYPpuTxQufM0f2q4d85HncR6emmUZX944xJmHsizAVAq2MDoj65HHC
jMRcEHO5z6nDqVSZW6MlOwLag6fWrooP5zysmOlTRFVcv4O86+2Qu0IaoXZkATUQuk4/hPwcMF6D
rNEZjHk10DtWZsOS/fj24vVVmenx2YDyxJi+3iOmg5y8HHvrmhx20iRetNpb4YmCH8mCOB7bCwPw
6n8vumoun6n5yXPejI4CokIDM8YLa678RIHvtArqsxWzI7WLLi7xI/iRuZw3Kq7o1o5DfCzmMemS
LXKFUTCmFstvjaviPrT6ap6COtZBYcEZ6Elmf/8n3wJtDVllIsMxTBWmnipGJBIdy4ti6la9zbRQ
khSz8rLG48e3SWmbUXKia99AF4SCqXhgFdHILpscOYL9/acF1RZaatmDTJlufNIKsg/evw3nwZtn
Ot37CGE5/h/c0TJBXP3eBX2O/RjNCj5Zz/nSrfp9rLH+D1FTZdXGX7+DtwwGlU2gTtApZddxNOMa
nferUJVOdECuFT2Npe5cu3OKrGDH3SbcW88ncaNiNRuUnZP9f2gn8c/v1nubjJEvVbUajl+V9o7v
DTuZuu717pgsvFdJMA+6z8E1FvgIDJpw/988V75OlP1Ed5H6ekfJGh5f8j6p1KIXbx6BIFsEJeUS
14m5KZ3lxL1KC3468oi351fmn7FIBJ5G9FaJK26Mg32etolthNP3Bwdc9Hb1+ZcMQkJbJ3iDr4zE
nwWxe4al71cSJoTJz8gyLWja4SnA3t8S9QG+a2OshlH6YDBOMDeFEgqFRS9FJpKfcK1W5umhiAyr
vSy20KtMdK2sgsYelkj1yD6dHw7woycpzBwDHEmT3R2ZKO82l7y8yTn8of0WBGm/iUB6d5fxnNhu
W6q2kIoFVP/sTIlU3rLUhlgMFWDCjLTCYxMXhilJVHyJz7amFTosaRJU76JlJmsHRkqoq50C6CBS
nQTISYNwalFGWI3LzhIq7iv0exLiPVtm2d7nSRAUylJ6ELyIULc6nFQD4RyNJnYKCstHPT4NZluo
wZM2+SXKjWI5l/BreCp9RXSFbX4VKlcntsDTxdgB+Pvp1h8DEwUVhuO0oabzb40PstXkk+krT7Mq
XWI4crGU7Y8xSiyIdu43tflYEDJyCKzaOk3x1w8rNhAcIrd1Y+88uK23DgNZsw0VXkSc2C2WGRvl
XY2PTXVdaCGTog8WyEegNOIMI9UoTmcWJEhJe9AA7URJp9DVezWu4uCWHLfOvwZI7qAyubmqBJnO
2JZLK4KNcIOjg4qEBaRsZHEg84uYahO1ueRJvTgRiQBqti3WeeeOUoMz9wYFRxA/1dsNMG45zKnp
49mN4Rm86vea5kQ28MTS3TPU8mJRT2Wo6JyrgJd+onGuIDpvpHIGdPtBkvoIv0Ecr2u60kXvAiLW
+n52sutBaqrcEIyuyMB3LeMSaGxs5K0ypxaofInwxc6natdf98ifDTKbuaqU+T043aRiLnYze77G
SIn8UfYZiQDA7MTrmKA1nOIEE8wAz8/zet5sHKCOHAxbcmLqX7mxHu86qpySKpH3vSUaRWYKn8Tm
mU+eWLZo/LQMErcBiKtgn0Yr068vuPHvhgLav2glloLANXIA4wV0Yv7u/IDHPhKtnCjy81VU/PiX
aujTx3zig6MXbZmir7OVTA0GP+5NsjnQB05lsQT3t8MOL83ZXICgEXlOaCHFt8jryUtxRuwG/Rem
tXVrMTNUKoM+buPqd/2JbEKLEi2etl+ir9tFikheq+6R1ccYUZYC4PWm62L0vzRZtJL0iH1N/8ZP
ZZ3RazbYbygljC6W0RR+S8gqQTVQ0IUs6aMrlKg+n2v0ffH8CAokywaJ9vjsckgbyqXfPmNZW+yP
umQUa7GnFGG2FdDDOmaHp0fnSqZ8d4vR4Q0aMUmPpq7NYDFHKcvWgftVIhqHovWecSgmlLeq5wnA
/XGMJCEo/PX/gMehkSgEf5Xmrglty5mkF62KpOsOa2shEotSziG9BF+9DIQ0mGIH39zXtHOif+ju
BsUUE4zNDR1ZKfKPVkdT7oU8QN7gDbyyqP0gcyPNDqXXpuIYLkNEiXOvAIx72at3DalAluDg5bmE
WOHdVIItWV3dXu7SeEBppb0yq2QWvlQcUMWsXLjPnWRMoUF+E5+igS0SBV0H50Bll84a23kDmMgj
ff/7Kw7a8yEvWPP1HopZBvFVS/7Z+7KFCCzEj2h0M60H9m/VMIKUAFeOY31KuOxtKoLfqzIVKBOv
Z4iUmZ/IgD+e1OBS6CC/TibyRMwhykALstbu6InctN2tBSJMg47kzaIhqr46A4hIPBgtZh6ImIWg
XNDAh0UcWhjk+WJWXBvn4l2KtobcfuhYtUSvqAfk79jPmyhfjn+j8CbFAtQ40GdVRKHQGPFdVIql
R5sq/d3iw8QeOXf3EqdBNcSJLrmsrI4w5mGYlKeN8e2YsPfl1OJkJDtNEX2RNgFNcEl6YbLXkod2
Gg7Ncy0ekut1l3u9+OmOcBTyHr9Eng3xlCaf0i/5QzX6vUeJAy9jYE/mQiXrGLlQRuriDztw5af2
oOXCOfc/W9Hsi9U42e/0+nAW05KqZShpX7GVrDUH0Y4/jy7v+klrs427MNTpA95ndqLOAjtNOPjd
9ayDGlCa1BiuSUkKGOaWraaMMSqGY+3442k52/7Zm1AQ6DFiKGtvyHEyhKNPiisrA9TAKserqrxs
ifW4VhLhLiW8rmOyJL8PWwnKMJGuHEZDy1/glXuHCT7r1i/KwvNMSpT2mP8Np8iFlJSZRfv/E1st
Kjf7Oxp0t00nx5ZT3vbDiMAUBialimLG3YAd17UaYRbWlwkzjlOUmabGihYeSeNt0nYJTOlpZ4uA
hc3tqNBN+YTPZI4tGf/PsnH1gxvq2IpV2HubtFKsYinBXn2WJY38zwRIrEvOuHOCBHE4/T48IV+R
wMmZm2lT+5LTqaaUSi//FUAmklZl9Ccx+4he/28DK7IXS5gqBdVwivMp3wMftNQAXC6vUCvGIK7j
SRTTwf2Jeot68XAQeVGgEMQSX8mZ2xuOnYJnUTWDvr7rXqpKCQCUsb3GRWapDcGvuNKLLeeSVnqU
INXWqpe8a5h2Pnxe/Ko9jQNif8VbKZLxZahETqc5y0lcL7P3N0R5+BX1kZippaOTfOATzoBiYzEc
KDqU6nK4tR4vX+BDax88BWT6/Fl+RwK+VdYwftlK2bwNxLMwE+GU1PTKTqq3ctAvXA1yqDZ31SGu
r38fEOsRT+fbOBsFLK3FMk0LFpO8/3aWWc0KoPk9PxR6GITEQSmenG4BZcTqLtZtomIbnuejOBrV
khXa8+RQr6vIO2KVH5bq6xl6zmzwKMONujh0/etK8MoU3h/gFujN8bTeeVlbzzHhmxRorQnnefm7
shsYvetypz5gOlFLAs4tRjHNH8uQv6JWPaHmpNivHwn1lMBUvFDjgXAU2mOFmGwbs2i6avLOdBDN
xq/z3x/VkSYtTAe8YUOOMBqRvXCJHRTfHU+waR+TKHAbZaDVEVBpmK7AtfvKOZZ14Rp2JA8QJtqH
ybM63dMW5IG8x/0ziWmqf8Fl0Z+30qG7kcQcokx/a4H9FTUd7JPVNZrKZyn4nQzxTOWi34u5xcCD
KKp0DgE9m+uBXCGT/x0xWrBwLRa/0GxrJHTkvIzXZzLw84BvpHL+Ej0ybSCXPO2DvFyZWhoIOM6m
24l/1NB++JcIaTK/98GriDkaYtW6+YVIO2RCy6Wg1zKKqgLkAAnLu7zXXRFANS8Ue3Rs9lcZxelW
LoT1FVd2LP0Ravw8Dfqa/N52BanrIGKCVh70+y5T/N3JP3P8clQ/YSse1x9yTgJ9WnQ0VmGCvkK1
Sp1DK5xkucmizIcwjBQA80rcaday7Iu/KFUNbDNy0viYpVicV4xEYNQRMJXR+STNh5H93HeUFJpi
FB0LZugWUWOio6fxBO1lqa+hcDoc0Jq47ZmBVEv5cVlGbmW7UGZyCZe69V2hFbetVNgxUSGh7pAP
1I6MADMVxb4uVK0xcLSnXy42sxmNnRdc4aoJtX1se0kyiGEr9ZMq5IVvkAUgbFqKdFEpmAASPBMy
7Gv1ZLSYH4C6YX0XEsdrlOhtEGMWoWxfXU2dZpSvfdIRtjeRq5qq7VJNygyhWa1DqMDOWd8pfMZV
uIAijTOQ4oMMIjvQePQnROkoqAHaXagJbUmmHYUCegDBoSGoT0OOrZjMG+YpmwuPf+n1X+MTrDut
msmMi2tKZbyEW1gNHLFNQveeh5fY+ir7amPwxPvTD0umFp60iDGLjeFYXggKLWl4gCxtv2r+zP0L
NzVmRV5YAsiEG4pZfEO4zU6SlPSg/7TcM8IZnSJrteBLrr1TxkW48eKa+8vhbqbPYJZKMA7tfbBl
aRzDimRnPOj97L3JBC15HenFFJQPthvpEqGYeCi9gtxs/UuWbvfTxa40UlG2NpeUkWwxCRAJrt0n
BZJXgDF1puRBXyzbQ3bRDefFdc6K7AA4pftaVLTN0h8wRjJXaYKpG78C0Hxi89CGB4eILujhuQO7
Sj/URe7w7fI5bsUD0VgYHs3JBMy+d3FurfWk9HsMOGwyO1BE/A54qlJU4fhMOUPu66DAYnEGUtEo
0g3KimH47MZtrZMt8TLCAeeyBrXzcs075463MoQKeYZZzfRoe/ApA6b8ohv5a6e00E9b6Cg90MwV
RmMJ10WDeJ1FoOijQVSf4Vv8LS0ryaOXEhM88vgbxLXhh1IFoEOfQCMsNqAFHoAlzzBg6K232b8w
rCN8VwX74n32y4+5uCCu7p2OTW0K68sRWWQHmw3J3m3A2P161YZxv/ckPcXiLiULSTxwlk/H4Knj
zKlgQgW+Jq3fzyetC2tSv7yfRzhTJfvy26BCvNZ5/YpjkMNtldS6pr+reYkH6l+korcc0gXwbvY5
V9tZ0gahfmn4aFRhpuS2bJqBWWzEEUZzljbba5+qlXO4uDibi7nnFSWf10Gv57nEmDmyHKX7YUKn
beBtITlMh/j5cprTss6DKfWmX9K5yKix5725N0diVvSQ+Qq0Qv+uTm/FPR2BmQjDuF7PU77m5lM2
ClUXQPeDAN0NrOxp4tlQmsJxxoAIzdmSx+kijzYydHFMXTnuD+UlnYW52vxUpgjNOEBU4Gy2JxyY
Tee5NG7J6RiTY1tnAEciEC7BywtC3VikZZO295w7bZYVdolJfVBQRIl5j8M1owQcT63nxy5x6dWA
bOjn8KOAayJjsSd1CFPOYbiGG+zuao/Ll1aNV6PReC0k+yu8fHwcccSr22aQfl0NzjG2na4RyPNO
3FrpYbGYacfJIhipb3kwUG0sYjD8K7P9PVkAI9RBEek8VKGyFb89wpHwmsoIZe5UA/aD/ixZs1lK
LGUSCoTKs7H/CONtNPfsshP8CoyV2yOrKtyNUsLF8rynr4IJr/VOxs0TqKAZyT2rc7YIpxmIbKWp
aFEyO6ebf0Q+SUxNPvWUOpFhzVSxpHt205EmV+A4naXVwjRhw+dnbF7AYIPyq18bplfd64qmmVVT
gfps8Qp36Rq+oL2SVEH5Fged1AyeJSu6SegHWRoqa7SfjHkC66XcPQRnagfp2VZZuQiOk2Sr1mXP
uEXMfIFv2g29TKZB4G4kTck8QiiVw1YOpon1/wUDA2iJFZRZJykfl/k0F3GZ0MS2Nwkow2P8RjJX
w0lLWPlksbs8Oxd/fC3xUvKVWaUfSlzOb3EL3lJxcqDkfPyn7Kjc2Jv+RTL+w0wcP624y0IqAwln
sHKxneflJHTav+MLOiGEpRMvrPZ9gKUMUDFUY0TcLz9LeNs5/Ge2jyPMSwfWJbYXcpcV0IlLxdsg
TGN4fPgzqGuGue0Sg86xlkDtLMPQpyIHnfIUmheLoBZPUwgWIT/4cBDAID7tWh4iWHeawQCae4lW
YL+jgvkBsqLD34eNSztx6lk2iI0c3eI1ygU8IFB5B4bTb0YHMzP75xHTdykFI6nLYMzIUjMe2Egx
M98QVmSqCY97MQ5hWih9nuvT8IKCcSowFQjNTt5UqtfGIy7U2nm8EXw1a2ZvlhRFL1P5Y4fVeHLf
WlbOtOzyLsm3VXLo69/DO1BOXDyvm8J6yeudFnyGZFFw2ytYYTaJOUnAT3EPphX8Na1IeXn76Sxt
NQhA//yQlAh8DPukA9KTUIrIotCOOzxqRLfnxIhV9gZD7eRkPoHFK7S1ado8npT+T3lrUPv5oReL
1/dRLYH4sa0wmLN3n58D/qvkILrdArNMcrpyuntPz/VSxCpbMrZPHQcrJb5T6pu+B9fp2z/pMATo
sDpEoQPmEcfpeMgFioqjmQZZ9GxfzhxVBjxBdG5Eteh917nrc+igjFJK3tFELvbvAm0P719lWrcP
AbyEH2W+or4hzaK7sHlbM+91+ZxMRRet5W+j5YEeVThUhDMIB7o0sIJ4cZwt2BSo6TjJa0d+5U8u
LV1jf6lECUwYIM1rdGDbeT0Dl2iBFA6OiGHs94dz1SjLtiWnGIt1xUymuryBdACMl+AnJcF6Og0R
AZ3dwnJzZbIxkhefv9EQrLddtuAw9i72plrpdiHbmJxlfbGd7/CrQV2Q4jAUW2KEBk70XqzqQCuj
xFjkhes6W3C1lNNyPkTCfejq3xBEnWAgavkPKMO/IA57jHDqmumS0hDh3YbSOYH89QbcEJYoqk78
4oaxilMEbqojPiM4YEJbulIc24CM5lS+yIKlNK4aPPWR03F6VHlCXaJ+xsEnILAVaCffsIbO2I9G
v5xydEMwraSoLpPJHS/sYajgiklo4IdNnV9muWPIXXyoSy+aBxXLiGqeNQ62on39B0qchD0FVPqs
Z54XPM8i8PuZd1bqsqOZ8FIEXwT62uHODKQSfcnf/QukINx3Ty3t+Gv5wB0htC0dv6v2cYge3Dq5
hOtg3/Y3ZZFgf0HqSd6e6NzjyFGlwoIaG6JbZ2aAmfGAPeKq8pQzsue7N2zCYqi1xGrCFK7Njllg
VtILoapqQTpMeKR1TIPt0JaCyqITfxkK7nkiG6vXwod7BfiW+XWvJSOnoUtu1RRNXm996CRYur4h
/QdAczZT+1nhltZ/rhyLMzF8ymcIneX1LCC43iUikpftDahBHNO95hBkE0UpXs0X48yb869YecLN
V3jjS25i7WH+kX/SI0zdLv8W+3u4cUZ2RuCVrSHVF+jor7o1XPDdwUdleK2yeyalTUG7CJxsGCe1
+AmbbtheJson3qQLqzZPn0ajzh7ZFdz3bmfbLPBYMZy0fkFKPiuaWXl9rywkjojXMPpRqn1Qksu5
zMaIjl+T1AhQXzgD+9ZFlGMovQ2bKy1Lps3lx6bVf8K21ZxD1P9AvaYoAoZXAwuorpoJ1gSD7v6T
iuR7H5rkc688LbRBoYaWKOl1Nut08iAKsAypWA+JAbACrbEkXnuE85YrRkTnqpNl3MVuwU0tcscF
5yhJ2T0bN5zx09xpGZ0Amf/Un3no4ieTzULbwzW2H3ogdcWncehuLFWbdGfyaMqOJYPJPF5cKuOD
9Ksv5xFfiiRmfMXZEXpN4M9iTfiRPIKJWTD0qz4Sx8KRyhKsBWaaPqh/B2//pSgiNNXAfxV2fE28
VqQinsTWq8EVLQYVxYewl8FtGFdTXuSwv7yE3HD8IfVodY92gx5e4wnJosUYrZ1zYdiCx7TZWxFZ
EO8DldIgCIIWXyU4j2GPhMGvdW+0MskZxHrTQzp+qmWVPP98rzZroy9FHguO9Wvj8RysthM7aSXm
xBDUM9YHs6Ah0HSZN0rNYPyN+UFZ3i6rfTv9KiyVbfDecPoDqFpGhlWvAJnt/I9taeQoF0B5bT1D
ti14Zo1/IsiOMyrsbvt4t1ohnqHrTy5/4bwhHXqLeQfGdQ8MKNejPWEv77pps6TF5kPllLmEKnLS
CmYSgTwE0ZL2AVMYxWUNmV8C/VN3AHtyKmE3HDrBc+epMO+ixcoGsfhAqHDnGnMOqnUdt9ZSNrO6
kXuKS/ApE736qwSW4OTiJzZTaXbKeOa2n6to2ve3aZpyaIUSJz7HQ7yV0Zd/54A1KjSnj8ljZZkh
KOPKqz1FaB7AinbsZugsyd0+0JqyS5ZNm07up8diQdOZ0CQYGkDNWV2T8un0v8bMCA7i6en/nfAQ
L9imaZgfzZ8llIJOIyHWBfxwG2nRrFS4fUScCfQApC6Bg3hTl3GgsdIdg2g6oDQCuKDStP0Umcut
i+WBk6D1H483s+Nf07KeY8n8tW5hJFW1nwjr8opSq27QaQDMcHOE1uE6lFFI71/4xxQx37pgn9xn
FRs2qV+UauzuRlSEmT9HIlwDU3XxvbtulUpJuZq8nlk1WGKBEUKGaftWDexg3+XatrBuBc8AvSgK
TFNskSag/fQ5v9IjpxthHlmFpIVnMvjMSKAFCVzIQRa1jQxjutXo7fUaLf+NOHN+5DXcGJIPKzyl
KBrxRm+OE7du55CK3i1OsniMmotHCKrYekWfyGiaVYJIP8Aw4rwesGWfBNM2/8hzBxntVF5PdTfX
6ACh8B4FaZRIIu0yQ51+jGQmlYgJ4o3QFJcjvv5KU8e77yFdWOUTdjR3xvCENdp2QsnhfkZEiNY1
zxcP+WKxg4MntnhDaJVhHcjdi1hJkAcOsqXiUGfQ2ptJREbGcaPouaxN4wzyK4UehAkA/evbPSra
nkRuVVMgks4CSktncJMMcc8yJUYHGfcM6lZqdHj5TAMJkrpuDqozbYYMgKbaZsuMbb2KhR58oQ4w
aQ5XoTD/oJurdT7mKwgo8GggtVRFoa8u1RSyfgw+mEu7BDI00/y4wMXf9jyFbHtLwg12U95ZXEaw
qGeruyZZ3LmlaIP54vmbsAXZxxh6Vj0yRZ1QDt7tj3VpPZWLLdhcod3LDFddIsIAas185t1+hFER
aNM3qbDlrt+4h3VerRko0W9E+g5Cci7uoUYurcdkPDjghUrnGVHeLfQFWhWqkO6kilV2P9rOPTRk
FOqb6HNdN5KvNkqVHciOILPr8LaxCPSZVf/nc1Fdwkz4hMAbtnTPKbHtiXWRNA13jHjDydEHwzED
ORrYi7tB9h3Ibo2+9UsY7vp6qbB4s7spdOuxCh4Mazhetpp8TDTXU/1/fJiKxuMEfdSCE1whdzx8
o4RgWPRd6h0BMSaX6MK/qUGP2wQxx4P2wfpIGbTrweNLKiYzEB7aBeT0epZhL2Q4vBT/1/l8LM/h
eMSsdAwn1WyfKO7AnmqlU1vi+FBDl/zzUbUHIwoO6tJAxAOwLd7m1i0V0HHYeLjfEysQXQ/z1WqS
r8+gVRCXDnPUw8T5eTw2QsWrEVPbNIQ6c1ukt28BmrndrwEOYot2qu3CaviaG1/kEOzJZ6qzUPsH
vjnugsT380E/kC9Rci2lsjQqmtQW4CE6j9uGxyVbZL3Um8f1JOmb4vLUnzeqfTNTSKaFh4zsJa/j
jL5yrO+uKix4Y6fxWkjo1RYn5ylnFuZ7FfwKA6AQhq13Ny+gFbaxk68RYF4cx0WgWnGbx2gz6u1F
ni3RaDI/PpMwxXe6u7aie1ro57vlCaEx5Gqz8ycfLZIVctcpoSrbiDNhpYMk0necyzSrnhwINJgD
4T5yTVuYsDETOal3Lq/oel7p5O/TUJzC1iP4Ei0lLXlIno/0I2ybXvKXDMvt1fwc6SKVEDMHFY5j
agYtjXWUalig6JGU/KRRKd+U6z4plGXFtOXs2MLTeFbvr01RCxAbB9OxdSppHZsGhe1uH4ofHLjV
+wDKuMrLQYSezz10k6XyRIXvsIfZgEZpnyy3a/5ah9zsiuVv2uO+bpuFtfTkrgZLDZ8ZFy96ISgd
32TALz2AVdwi14jhgzc0J8yfqYx10hC99nSIFGL3yGDEi8xSHdu/YicYBUJpgPlHUJj/smvnRgVy
sixHLjprgLsK/DahPiDrHMppjEYdxLaI6yZBrL6HHOXKZp3Nu7U8B9XGZpXQzDH7ARwqeLZPxRTT
wvhpiFmhQMAbcCbrNOgy/IxWCm7pxu1AJH88PxjbS3GLQ2V82HfNIbsYKfNcJGJwrM6XBOxDs8il
xDLCYbe48/ZPX25VZEr67kYI1s28ESYmDnF/EDdxZg0BZ09ketBfJKOpLpIRlilA2LrwuvrdaF8v
FZ9hJje2nfvMfXxf6QiCyJ/S/SW/kQkSqoMLgzz3rISDEFOc3FIwAxkbhBrbl4uOtl3rPcsEbQvP
Fg0Lun0+R6pQ1xqlnwNKB7lmuJ2bYSz8WWbx/8nE5CEnWEosXDOzUD6WwYgBPL2OEX9Qj7teC8ld
fgkrQZJ7sycyh+eaRq9c/FFPNgXzHRxFU3bFBz40skJ608Yc5t8hTcBBYH8jmD93nmV17GuRxYsQ
nZ6iq5ov5PSp7KyoREszUi3hOQy5Y2tipJEsaZgGrJSWxCQM6fGSVzGMulpaCLUpJ1s4RxJRC+4P
OwUIcjc0oGeFLMgGg7YzEXlUiXcS9lIK6FgXStqzOgHSeezFhsxhAagBPQDFSjLY/8xmoCWGU7Ct
2fmEf20jQi6zJoH/KS/EmXzd2rZgNCHP2zVpq26KdiTBioLd7Z8/c6kZKqLWOMFYSHWQWCKnVb8N
X3QS8alby12yj45Em+ZKbTNPjJMSM69Aksz9RHHBAHIgZtp+WwAko8d5E/DuFoQnS8GkIQD1QSFt
MKWDwroQJ2+htoFKyqIgtuwOGS+A5IUVMGW2N52+tRu7OY6eBufef9YUAGC2pqeeZFOmp8IUUMu7
EaESpwQmsdRIXmNk4zNF5D1h3NXgxwfXZlqG31fA6BdjPqQL83rjQAiirsHyXF2nuOAPT7bHOB/1
+H5nQA45kXyEUZ37MUJUqVCk3J5GNZiOyp1yo4sa7jjG2Zgrp6UnsreVqVbBrFz/ykGhEbg+3bY+
RkQdq3BjYJXJlthB+vSDsZcqzdE7Fk7lULuP6VJ0FecB/+kR03umSdmOqjIEgDjSD82n6rIDdyIM
rZ3o2laaVTo/QBJ94eRqt65tcx8XN+ebojpC86Wk46zHWwQQfNkivZVbi5sXCSVrgIsM/Rl5VLdv
y2Eh93CgsNiDMYM8nWcCrRTkx2PYWho9vdixbKLjrKx7xp9y5oiW/QkB+74F//cJZHL+tHRftnn+
effwghBOfbgVpKZzfpi2z0Z2iu3irKG1B5qYbvyTwLlHj+c2UDZs8q61/UI9UPDkKL0tLvg96R1B
Ad/7afINs65HuDZ/1VZdBmh3RT9DmUgr4Kcevb6PYrI8CGA/BF1bqjihIXRDbbIQyQt4BllGjsl9
ttsYkE1nNmq1HHqx1f3JTwsrcFi4CNKDW8RAKoEERiBFrc1tqjZ5aQdAYnIqOefHDurBq4km713f
uKB12B/84lowNI9yvAcbVARkBYQ0U8jzzluEmC5jf7rX+hBxisNyrITvsHtKiSFShlrXsTrxLqnA
ak08Gm0EtJePQoPiI5p6kzZhkOM/qBFI1a2HyGnlPX+b4CYIS+T9EaRsP0/2knw4L1hZDGyLpqCb
LoYIV8BXSpt6ll84IwaERC00xH2rG31upwELa04uzcOldkCEU9R/dIfxysLHySg/B0W4maRyAGcJ
mGcUNaa/9q+8WqtsnCwv+n/x5iI7h0xXidqcpmgzMNfjWtbWpWOJomrCldoJn2Y7UsqGl0sIsGnF
QfO7O8a9xJ6smzn/lnj9fSe3uHh7uOx+CMdzq4KIghZ0HnS+QLosCRdWYmQWkbeA2Cv9l1fMQuUU
vRIb2aJGfESq7TzGXqoN3Wkrr9MVJX1SQjPCCuQsY6wBI4fqu5IabIJiIlgw4XFKpgxZovmuF/q3
ivYawyRHCHB+Jkl3Ryeg5U7scdBE96KImiPthfDeuX5kP9ykvvaToSU3N3BFbADwHYCtHlqATte1
2AaY4jAm+cJUMaEe8aT8Vvqy6Zr7Uajnago5M1fWWlxpbsoHVjUGTDxRYpPG+hdja9f5+K4HhKkx
mVXKY9bFNp4HPI9xjkY+HNCMe/uS9+XdAf2gNxKDXGTP9FHyVgb4JO7j45Vnz1KdfpLvDkEzGfL9
HqTPe6M619MI5cWoQkytiUjIKCnQnJ96jNA5gXq8ldMzn03M4+IiTgl1+7J3/wETbqzk5m5j9fPN
Q3LfajwQfCUekGW19MAb93/K59NQ68oh8f4NgpLlaQQ/C/dpx2lhOGXu+P/QDXUPSvIYCcWFFYUf
EXbfliIK4q8x8JrVsFXGI9VdOMZYOaeZQ4LA+qbwjIaCNBHVHvriqDilruWqYJouHIBXc83QRzQj
Bn8WWcbX+LcOQIQceTosW4GSd1qfOp0Nd5IC+HhyZafYohKV0GMV67fpICjOHA6GbuNsBM4eU93a
mheKJ/svqCMwUgdnfaDVXGah+g5UiWPypRXpk79VHQqg4ecG9wwi7unHXcQOz0s9UulNohPknuE8
m1+2+PK2EPnbXGQOSjOoQ+IWjC0gvxQH3D/R9UAl5Pu0Uudj4PQWJ7gnTY7x2IWHITcprB039B0W
q56cqVMlRz6WYiUai7cNeA3QOhepAqaac7V9ym/6qMXMQ3NLqNqPwLT3el5eme09RkRNTAdiJ3yb
nnwfE4gPABVBZWPEg2dpF23UXxpOE/RnGzQTN1VdorRq5kxogjQCOwJNjeOZwlXUxcfHyHFGT3UU
RoMY8d3VKSPeNZw2FPh6UNque0HeFfUBo2/ERktSDt2PO94qruqNnfMIMg0xx9DSWCV0XInYr+De
uipU7pbgIg/RrkvwegZPgnxeAeA9T8rNRuVCK3a7THZvvrQV3xBj1Ip37UyYBBAu/xVP3Nl99s4o
qo12vyrPoZmbiT1wsI/OT2iG+ShJA5ZXh7Gt0uIAJdJTtFx5if3FOuFQh5IbnWawZa8qCnyHmf7f
CYXaYo1Nabzbguyx/UQgvSqYLXwAeQiScjiGaxKjykq62N7dkYru1Ckqjuwlu9QvmfwBulp3v2+a
IosxjIC2BSy6uX5zDa9E8V/R1WFHztyZPB4vpfsrXabXbiYTiVCA1UpoClExTKxAwBnSlZjFQvEr
ICKIW+V57ERdSf9rb4NbqCEs7kEs3aG/nN+ie6GoN5PfnjeFW5tnBgdXDHAVRsLguN2F1RuY6CKM
9Sh7ZZfCNUbp7oh1Qfld4hDLQMekvRcL3MlAzSrfVa3/MZBgfE5sFP7+oku2f96B1scrxylA+Bqv
ZYrSZA0CE5MUK4UkP/0GLoAqLRFFVEosfIeuvs3/RyisQMvdjo1Ogt5v0zR+hQ4Pe7q4UkRN6kiD
wplDDixihYbgN/7i0sBhULWeuCq8xnL2AMFRL/+Z+5+b2sTFTLt4ntmtmvVzB0oX9VtJ3HKDs977
gjyAqzkHvfn6gtkvTEdeXwnDyIb53Q4r7gkyJS4L0KeFD1dFYUofCCL33IwAaU0x/MVqcMx4Gpm5
bYsU7uDWbEJ/sganD///qMrp0bIqQOQDYW1SHLtA1dpROI4/4gemvr8LBWTJC48oByE/yN1kiJJM
iYrcrFs3C8qyqRMFq/6uRXsXX4ns451Ch80jYZDqqc3fXmlRFQcfooTWhmtnsD7WQrMci1vfi19c
s+sa3LrDYIbhbIXqq3EBmccU5G9gEOt0tnhfLZSzmLqlv/jbXYu7oWu7iU5NPQFHU49O6j4aVISb
JpMFFk4Fmanskr46SquABoRGmBXNbLVn0Kr908If9OsLSoPaUcMXn7ZhL0yyBtcIrU3951vlHJem
7DXZC6ymQURSMTM36l94DT6s9J7P96TIYwZhD9S7BsLf8fZqTSTqFUXTLST+Xu2gYpcTLvx0tIt/
Y9maUDhZ5l9LpzgkchJjS7f/NQl953qzFwGuVtb3tq/fsqbA6jxK8xVALnCi6mGnYTBvEAfS8Uri
qUeNBMesLG9mt8fpJM0vfAAifoRZ4qXTvVZ1wqIId9rKbe14y7fv+S3dI8JxvPz6Ky/Y6jgWXwf0
744xzZg3AsufNVM5igePcRyotETo0WEDufn47cdqudXB6xA9/R45z+j5KoeCEI3gjqSxdj9gcwdq
h2/6YFbmY7FiYq1mPm7qsKyNFvx5YYzoMOwoI0+W9Ny4diboGuuuVhvvUKF7ObEEQ2XIvS8hXPf2
fdNpfkF877jjsBburRYpNOvGvjP80QUFKNxs3+TnuUXgs2aYld2fcZ5Tvl6hVQiz4H4C3AXtgAUF
nLodFi5GKD1eorwfafpH61H6RAcYRAmgzlJMVMDzGhZPpQJMxlOU7lXAm7Pb3QTP+FBYmkCpqjAl
m6+PuCkRcsadY+LR6jxdtL2SByh2PPwnZH+X7NbvNox52OWzS5W+K80MQSC44HjCyGoovY3KOSyZ
n1DaclQ4tL/p+NpYtTZh5SJAj0LFvPOr14WJtWpIwpyqePUk7JI6jGKDpE+mew7eGDpRpOPOuvPO
0fqTutg5b0SQHIAqiHd83ShbfZNarx6tq32F15h92kpFvBpYgvouzfnNTXfHbFbzd9Kgrm0PoUnQ
YN7M9wN318CQAbB2pDrI7zs9bob2yvJmbGOzzgquU8EVKWoqwRu1PtePRQifY5QxdIuvyDB76A8k
psJQXfYh9INmY6aUWfYT8a11r5EXupd+AShJ7xsVABoXpMuFP0ybESnG/p3P1NB7Xiq1uig3kDmO
jtn7BBXrUrhCdxexqStGpUmcLPg8ozPf+jrWL6wRD8bWRs+jPkA60ExQ/r14nRRmduaSrMm+GXsP
QN8i3qdkUDhBXCnC+rKRw3kZGQgH7RvNBXhOxoWs3NSYFzK47vXGepHvWYVHwFqWVujSxOD9/JLS
bxlg6dFqMtMFzbpg9DSR9IMDTj/WDY/K/qelAhzKVMa+GscvojbBydJ8NzoDXJSHAEuDNpk46CvF
70L+vwsSVBPYzimfxgV3baY0Du1ab4xBjShJ+GquPXSQbUJxynNOAzMQxcuXntuYdjsSWmLPTTFJ
GjP6w4qE5xiMetEyz/YqYyU536r8OM4t++3cilQVB07VZRSIUpGHLKj98qHYCa3S3TeXp2S0yZq8
/CiNRsSTrszig1UaN7GTwgvPxU5sM8cgHAKoANT/OmfnbsuDp/2oJciOW9Xnp9v8jBsn6qyGnWp/
mORbxUB+CXDueAQDPsXQF9eI59k+12neqVHuJS7Yij4k8HuZxOl2GQWk+3ILsVyp4GVSHL+ivijM
1XdxNQnJmNATzcV4vAuxRCCbhyXGBPfPCL3tRCMDuYcUK+YxA12GYsgwfM5fW7mj9L0iaAKlGICu
0X6NN0o7H5TsTfCV99DqpyZtsfj8R+YYvLNsQdnCbx8lzIKaOvSiKXWmLHYIikglLslB2cfp+gSI
RXsfl2a+oCYetPuHAWk9HNGHMW92s6m7uO2tRKHlD0E7IfnNqY+HFAipfLVaPyIlSvMtv1VvXOzI
LCqWdIj2sNRvxogZREF4PHBZTZFwVFFNVkQ6+vMDlkCUn3LMzha6cOAuJzyyBuhFbh3SI0SSN2kN
9jdI3r/GL2xmQUtBl5Eqy9xwOHa4Gz9CsmLbWnECS/1IiSo++z1XtochvszSWI3wPBf29/4YKbe8
Qs75lrWdlsC5ThsvRxG23qAniwTRXzhtpwLIVBlUHgaLtoyq51cvEmt1gv2zYc8qh6yO74mTx/VH
vnWC8wrugUahKSvX//EHhygr/UYhoysHhR6gHXgvB60lnQ2GqQpI5ktcaJG9fbZC+6WXtGdr6b2Y
E1m3Bz9/VK0oB6Td75BpSYSZeD5Jzf0xvp21MSOqRdY0DlhSpjaIB9bWJ/e3xA8g52vT0XScjmMk
KwuV1gYlfjOiIIkSPJDox9/YyHF25VrzWtwAajK2g2ulF/VSXa2/upayk9M9yR3M+CXK0LPfh4Hg
oT0EQ38H9Qzwgz/mwPuddBX4QC17l9kfIZaYxwIBOl8yP2s/oh2w3W3XbQMY7heK6tOTvJGQ5iXh
Zh3oD4PPBEpjHF4xj0B6u12lc6trIhhgtaABRM8DZQS6vmVrFHB2wmF9oq3RIkQHGguAcDsoIX1q
E+YEC5on99VIcrt1kn3fSBq3epSjQLISR5nTsmdeuYxntNE0fSM5EWUfD46AY0cSZnDM3uTu26+6
puYQK73d3RXKotWOPjqzbFh6OMfj3WpTWYHjnhwU4AYwcvHyWXYDryW478WqXrYHB5v7akO1t2/n
MR7mbbGaySmoBK6he5mn3bivw6nLyW3LyiAk8ePRJGszQAwIXaA8ff+SMO/hxELJFM4yFeH5eYLt
4Cb121GQZkN+2G5wwrPj8oGF2afJ4l54/Sc6Ft73x7X/dQBSVGlC1t1+t+5gXdxWJoeqRMNSdL+0
JkdAYA9iFD+pCwe0AU3iJygeMmDeMfHdk0rAjzbxt2tnp96qM1l8Epo2uMqFmCLc6iC1DcqUPVGd
8I75b1uV3v5BvaPR4j0qL05Qlc3k6P2L14IHqzEVTOGXiGmvq245z8k0CFrWfxdcUQpf56gdVwEP
xhXT8mokysDxrPgikvAHcFMoF2txJ3P7T7ZRTcy5m/hEUcJul0UqyLEFkC+vRaiaNIkkYdKGx01V
DbtHyiV6pe03hLw5hmkeg6XYjEkg1qUwzW13y20NT2y1Zig7u9jXd2Wxb9XGI7GRnqqMOTDx4TF+
8tOWMhWmFeZR8wvqwywQv49oYFgvKP4V0eZo/Y3yj0Db0ZifEebB2gIcFIezn3u2ijKSgDqhcAyi
G1QMCUjCHIMh8zsklwRJW7I1kn2DwvzsshGPmCUa9fSa3lCxX8Y2ZKRt/JjPouEsOZbDzNSzCoDb
zRLH74B6TpLuRKLtJsUcY2Vjy3VY9pnMbJBWl++2zemnIG/Ei8wRyYXPc9Yk318hHLxKIWzeSFfj
h6+nqN9N6jyCnN+2Q2wppGylJ/P1FQTbT5aSlFW6WHMrDttzevaiFxL84CmkOqJ4hTE1FHH9tnc1
ufPXNOo+EBw6R1z0xeOka1VL8PbON3qVGQZ9uZRe+XBUdRMZqVhUmuG5HQ9e9AKgiZtJvm20vZbl
HoBncdmBSohLlivrbDgN50kr1cw9xppwcW8fJf8llEFN3DMhUc2AJHCuVeWTYIrilUabfISohuf1
So9BCTRWlYYU0R+1+64hmPEgxCSficRxhMNegoqbRQeImo5t+39rr/XRfcQ+Gg3ix6cM+3w/ZQKK
L+91irEji+Q4EZ+Rc4c5CmqIvjRqqz4VaIUH38Qpd4idm7J4Kmuz6kF7lDpGCKq+/mzyzMlwLRsC
d6UxQHcq1Ap3NUmQghB/N5lOYnkGrOHpuPxdeIM1HfmXVcA0Vr8qmm3kxgRNW8U69B0vhlZPrK+z
qX36jzqRFdJpngHP6NirzMXnQtb6pWC0JfuWKpRMGk/Zn2n8Hc4dYJ1qsvyUS/5kruYVQMIh99RH
QBfKWav81DTYOUKAdOZL8YrtX8ukcUD8uU0RKr0Z0Oy6GhCp0eeoZW7RezIemplpkIqRwOXFvqZY
281TN2LavvqRls6S47Vk1kg4OxS9tF9BTMRhJNIllhqXYxJEZC/+z6+BCmlg4GxwhQP6GccMa0Qq
MrFecbBsXGyO0TRI9YxDfAVUmXxzBwWtMdbDp1Pzny2nMrvH37UWujtNuc3k+nfUGly2ieEdVYnt
dduXcRPWuNkdIzxKDkfBzUg0o+vB07+MbyuobSYNVwZE/FD+35MDNMWSThZ9bA94Dob8DGzJH339
gWo67ACSdZ2gVWh3zvfydoDCAa+xR4l3wU5ywOj9HY5i71MJS6nI/xwD7LNAiCzcC03EZ9pm/Tfe
uLPV/FIn+BWoKVs0zw3LSRQ7LdijerKxf9Hdwqb6UiJP4w6j9yGYRIk54MOmpgCzvQApse/Xb8/4
5ZZtA0oz3DU7KB/ggG9rkOEkGxnfdDSqnRRh8mqLuh5EzUFrc2D5Y1dl0gnUCnYSv5+eviMGXnvo
RJm8q064/M7Lo0XrfM/nB0TjShk5gWx8JTvEpQ2/W4gfisjnFLClo4rqif4+nuzgcofJLrnoglG8
/+45DuSfXekAeSfCyCuuRe29hHGD6RJm7YIkOlkSO4fyhhSLzsoCi13KFTy7FpViTE4LnG4N6H/P
S4FGn62B0Mq8xueVw+MHirJrdrgbDuKtVOfpSRk1Qw4gtINfW4VonlWeYBC4nqwVRHkHuMUWDyw8
ozCw94P3ZSZ5Y8ZHMhYSNBYa7hhxpWYNrDfTw4/kDzsaMyBGxssxwMvU3njfQ2D03z+Uj6liVxq2
sRu9sklsPk78u3s2nCCHNt25NOlKOycRswxEl9sTthR0Z5fAWxtvOmt1SUyEnV2X6i/Ll5GAJVRR
ZRHqwrxSlnZFeN/LCCCV2nYyntOxNtL9Ba4s8V1kLDfiS39FgpFjt1890IK12GCIT3wMwVuX5Vhz
5io+Aq7eQZXlN5t1TmjtxYpKjJ0zVMl7W2y9n7q0fAcpmeeVHlx11nSiKOsrVTZj8tpO/DJ23lXq
VtCedY3KG3YjqPwxpwOs69aks9mA2WX4GZHCbSfrZvDRswvCWhs29+NjEWgbQDUqKEm9AzRalA4R
QniDzhmIVXv+OeOkW/Q+jbbmU34gCpfDX6qPhwUpWAN7GK3vZtYo5JpGvenEn8LMmT+6xKPTOTRf
bjraMa/unfuVoCP+39rzz6NAUBVRFScUMVcyOcQophCf/rRrMC7FDbZI0YKFn0p//JdkTEJWbeRj
FlH/zUDZE3I7N6lLlVIrnXkQtfqtw+ZAH97rB3h751TwNDnyNLr/p3TMX20hFsI7YXZglSLQcnw3
XD5F61fR2xtpt/gqe7uFfGMaWWx/W5KypE5BMbBfnDMQR8lYzLzlmSeUBewAHOoQU6Zsckoa29yR
POPzbZd9gNcdZgYr+S+t2Sx3Uq/+82rK7AJ4DGOOPNqz22k9oL6cBu1qRhFH00Nw1t36Y3vfy5vC
vSOCiCDkw/nrWkAQCroJziUPOObiCXU9gKk3mZ1f5OZlJ620kkZwcdDHK7tTG5gwOmmj5N7RCtYM
JUEvesYdnw/3jEFoO46TfwCsng8e+jwxvJdK1akgFa2NCMoZm4eyFZeik7NamSb+B/bC8WvIRCVU
N3Bu675QMcb7BQIcd0E2kmtT6gryDVfo5Bo4v27uXVTU0RKOTOUAomSQLZJxZ+OSSafVrBnZv4+O
l7rfjbq3JkYs58oJCFOTs+dXFjo0As8b4QNS4usgOGv+oor9w66ZGWs/avkfHJBXAyMtmTOO0UcP
7tLKBTCwkOxRRpCscjiy7XA2n16LiTICuJOtbnC+KSuKhG/F9cyIjd7iIBHi2okSHcxIyRchzvOh
IFLp38j3pO2kbdThD4Zy5F5zIw5asadLBJSiWV81wPkxpYL0M7yZleNSp/ggZG21MEdgDyfVwuej
v2kuiTIs8UKzpgjnH0qJw4qIMrvXxN6EmiL8hH2ZflOMYMu3nGROGUrHbkFhLke/SIJBjm5fBTQv
zDVe5SEx0dc0ARjUfKGQRGOsANnNje6lMJoyk+Dz1G6EMqz5eOu06N3fcPNGICKZc/+mlGwE2rgt
6oBJy/Zv9Wg06RWrHW7ZAqbkNgDWts3umxjqwDQeIZHxDV68pCNzj3n/+wRpG1Z/WhqzFVtNAGVl
lY5iRNs5SSUtN9i/QI+H42QBok9fh1lzr9CZLbX/1QNUpQxegxcXbtjI6yK94ljFyI7OvC/RWmE8
Cfx4lXsyLwSJ1hiZNp7wp0jxkdC0qow2+tE+zXgf5NnxY0O+zrfEMAz88kwHfPWc239FmLrVN2BN
+W5+V0zpdeKLyiOCdgU5ZGPVvr2MUiFFN/UPbx9mEzL9zNkRl9fCiI/gvjExOwUqcQ5y/I3lz35s
hNTiCCCwJwB7B/Vi4mX7Dr4eOBhgJ2RTecff7jdKdVJFzVg53hWSRS7pKQN5wPEDSXpErAKZWlNH
6XAJ3OAut0SwwB7PlV9NKiJwfcNHnQ9b/3e9rToCLl7FKQLsPslAxo+ISs1kjqNftVtEWicDmqDw
FBnH8CS0ymH9KTy41bOqxlgM86hulewIul7i/tiWXXEqkiV0YrMsCx8e70br5UMGdJrxaZ7d9XAJ
MiiBoIn0I/KrAwrWOIgXaG4irHWtuHCqBaY59st1MLFPNmnI+3uh2Sgt3HXMH13wQogm/+mWwcJr
TiHIZV/TDz87vwfdpjj5bRwtEWFTY5IAXj6sfzJ+xmvTzNrv+4TQHYjpJYNxKdLgbg/k4y97x6lW
wsgFuJmAeipkdefybEGAaOBMW0ePiy55Cg/ntc7gc7K3EZ6O33NpNn2VwIWaS4/QaHrTabyf8r7j
eJhoSZ+x5QYzbATqR1Fn4hxj1hprpeyQtA4HHLAD8a8eO57p0yo+poXtwcIHcTuLE9I2vTVAF72h
vuAGFhlgX5nR3gat+w+8txZ5Hy2TxvnltQkExFE2j1W2IrtHGEvUivlYshJLpg07zgFn08LWASc6
HAFCiSAkqr9WFE2KtalzZWuRol8PljC5+M3RkZ/HSXEIGfViLyEoev5psVFjgN0ib4HJvHkBkAU+
jy6jLltYbMFz+yTZ1MGgkxJZCq0vEMtmBbMWvdD3cfeXoQj8Elk13Wm6Ia6WT4nfAGvtY8ffGWk5
P0k10JVTAMHoZBuQEnbP2Zzk87f+4gbjhmx3gAwTDETq/bD3yvvBmN94L0Rk95n1Cogtiy0ZE2r2
3mVRkzu+KhAcjOSPq3a/ciPx+CRQRF7aioFCEEg4/NHBbq6FgVu4CFONNtBJgMpZDetuNpSiu+u4
1URflk9C8dEwAaWFA3vGj0tj4IQR1FjBsQk5Bx3++qClML13ErzOx7CJecZ7U7DiTObRA0aF8rMf
+Eu5/mqn8crP89wPuh0ZaMng1ag1gDgS1dCQuDxxqqHBfp9t6OlmJPMiIuXyal94nYkuW8hcVOa/
zhKDz+Kb9BkCkxcJp/jvuFwcES2SIWNrjlXikxkQy7eRvodQa+mEvljTsy55LonmZ6aBwdVclcLQ
qkL5EA/lcGzCb+fdxvAmkZvnZ9bXWV6Wji7GBtzYz9t5td/A0cG8grm5ilOTqTAhwiVpwnNYDD36
+5HqFri5ZvHwWWTBwS2sp6C3eT1y+fkCpyfD5OOcVexu3Xs1KycK5g6ZOB+fhGVyP7TVwNLghMar
bpa7UG/lvxc9Rn1JCJvvBBv0EfhaNSuS3/T0Rdv/V+Y4X/d1sMVbBBKJy4BDNsOmmJD9m8SyER7f
TCr5/r/RRuL/VyVvihDlkaQrikBTLEyaF61gGC7NVfX5EDvzZPabyge15CroC/CNmuUTASKVp4N4
yxseaaZbWV8SkPydLtG0/a4KkvOOq5DDxMbLq8x51sLfi2nTnPUgc5aILJOvQEz4T7Vl8itqNjPd
j50jDu6HKDAEcq1TKMxLkiz/mvX4sQei40sKrDWDhC3I8q3VVwwCkNE0OnFyneECp2yq27SD9mpk
+ehki1S+V7erRqMEX13b46vZPhf1XnhZiN8pir/SbDvQkwK6dNRdw7/5JV3q5lgTorjol6Y8g15S
NeshEixgra+jQsgJrUCQap1/RSNTJD3S47pwGJsC8lTqoWpzEey/hIFb+3r0ZHlYpYtOo0vHkPUs
op0r7g7Lz+aPqmJVKBfycPzkeIabsS0hOtTDQq6n38C8sl1S24Wn4Z6hLMf+QRbZJU/Vk6ecG8kN
OuNWWBc6z+fY0YoAwe+dpk5XTKsWKPXUySXJebca708pQ8kxLko6RtCCO18Dut8AtXQv2pOwAKgn
p1KUEgmmt7OXnhepSiF/BqGX4415kgtALxj8GDKFN3a/KWT/tdKoGeDzIxts2XNWHL1abmQ2DBU2
T6PnzC3nwXTVYqo5uY00JpkvyQxLB3/cIetkPqecmUlwDOHeuYlYU59b+4C+3hwzBsM8BojunLFA
AdYE/dYiLzqfn/SKwzH9Bz73gKUIuQnsL+Hkzt6yBR6fAOfJly0LrJjGEpDBgnRQ+H6UUE4LEoVj
2qQLnHfFeRYuO4CrWRxa6NKZ8/pwLbXGQ/jRINEDSR7Zx2VT8IuHsIb8nIMEz7RP2VXG4iq9R206
sZL3xbWmhzrsNpXtCtjVqb9ACHQVunTz3WHkoqj7AhE9OECcQku8dHoPVonzj4fbt1b7H34xsqSw
vt4cgKMrCStFT+QLh/pv9iX7xf79SqDVK2T0MJvfvLd8tZtslM9Yst/UHQUscyiuaeaXWSprUBGk
AoJc+Lhh18yckUhczvG8qx2wAHmHMg1IbuhDvXvWc/QxEjmM/FjkgYZUG1e9A4WTuQ0jIqLFDo1s
fSHFmdwEtzscMiTjYWheqQAtP1BoRysQ4idvkCpcCMo1caQqBXQg0H6rsZgcuXvQhwW1vzZLRhKb
1zQv90YDo9y+dLrv4atqYX2VG2wjfaulCexKgj5tpfIQUgrrlEOxqyNx2urU9/nxZo4zoI8tW54X
9VKJvx3BnYxdFwxi4EbPF8QemkuDucDUPiLv4l7WI8SMrraHHlQCWaFm6kiAK4JiB1/wwVzmdZHi
iirM6YrJL6OE2Zu+ZMK9vreZ9L1UeiQpXDoBiR8tGKXJmsKzEo+U+yTWNOjNCwK1GEfDsxC6liJb
YteqN9oakfi7yNBQTYQOMjZDUr8p+eKP46qY/Pihd++/fTNpDVHsnMfFdQWw3P62TLDJJ/EzuOR+
aKchlAmqNUSsJL2ZUS5iOf7x4Qxud5Lddg8LrDH20WyCrz3fFv/LYusFIJIUIpF2xpk6eqT15rAn
NARDiF4JUH7bug+xhK/tbu6AtXY2qCYuyByf+X8wozs855NaPB6B0jUE97wgyz9GM5dNpHRJkKi4
uw0gqFwMNlmqj5hFkFvlQypys3eJwkieNPVhco8SPl3kO5D5rM4A1eNId+1VsexscivelSw7Rkno
ezf54Lm8RVu9Jc2w61rGdOexUciYGJI8B6t7xb0poWU9EV/GoHeOVR/cp+PZQoAyzYIbUTjkv9AY
7fVPrYmU6MJnP3rvhyyk0bROfPHbaj25prDXKOVlYqx6+HcKZ73CIIYC0pxF15i9IPy2Cx9Ju2LW
SIQpAIaFw+oay2BrJq1j0u5DTFu5RFyhM8ed7wdF9BdYa7rO/cWbn6NkVcD5cTecfEA3Ea/fJrvl
p/m/zUZbkwklLi1N545thSxFUwCT4aj3sdi16E6eHQMdBH2r4op70BM+gcbvUxd78BwUl9vnewc6
nTO6urFZ4KohTkZMreS6ACviS+pF7pSujfCkJHqB2ngBk4AMfqEkImjmCsNmL823zdNbq3qEbbxm
9nPK55cseIRGeXESVQyKyKD4GnY+diXWnCnhfoKuDcy5qPL1BGnQKSAM4m/Z95SDo3TEmvm/AVFi
DYjWY+bg/FKPElQX0mx9IaMoV8zlq+iBF6JukFAV/EWHc5oW14hiEqYU6bI2kM5ASRseTdnTcDHN
qKOxZ7xw/nXeCtHr3GCWrVvN/TsPSXFv61gjQ6V8FZQQDVqRWMlmOwWg4tQ683tky7xAgSp/P8ed
ULcoA0yX2YTHl88Zep+4KWmIgnG/AYqYffyqFp4ek9sQTSORjk06041MOSyvLx79YCRPQo/+VRcy
ZxS8WisM6V4umhN3w/wvVVBS1oBGgjQLq5QCYDMfGRFcM7yEwqr0bmqOdnyPCEHYxO+5v70xuZmC
ByrPqWUYaDWQRvttVh64Hr9oiEIWEPCBB35Nx90ozl+NhIhhpu0hJmwvlj7xCSg31S+G+ejBsEZb
x5Bynu0aAn2sFfjpAXaUrM28tap1AW/pqDbPmXLyvwzXXnOS3WuzylA+c/0iUjjqd5I4GyQ6tpTL
4auu1grdqrz3lpSxA65XzfBse0yDicBUZcpArPFVW8KNxteFn2HbBF24es0+uXUS9eqmVADfDaOg
GuVE7/8GLlqiHDaC4RIcl6lfq4s3Eriw+6KGegbue25ISIgkFZkqhn/9dJJ1R1cnAhJFDXgMjFFi
xlDDJ3weaFR6wMpKy30qpcMNF8BsH/ZD8wQkMNZLjbhga8Ynz/zXfptDz26ksCbzcwQvRCELTHAl
5tOvqp6qjTF93kxikIjw8t6F3qe2ty6Zg3YZdSjcCyQyUYQcYytr/Yns4uVKXGqJBFx3bJ1GxlTt
grZZXf/+3YpnZVPUvmn/F9GnsYDp8JxOnZUwOpI5awn22J0HleV9xTTa1KhN8QPekZQcmYtpjSWu
mMWaP2FgOhHPW+N+q6bFj+z7p11/bV1YIIObYwTmqkt2ZbjQIM/HUUfQsm+XbKcHlhjLn2pl+PaY
nDNvCduyEP3qEYsHmuTwKXTXtPDNMm5WUwQRSobmFX7GMhXEDCrmXnVztBg40yU9j049IfQAMo4e
3PjUY/iyuoSxi81HNIWq5pgqgOFtN0yWjfERUqJKuFmHIXDQ1xtT7UeEl1ATDOzAkv22iWOhPB7t
7dBp8IKegBS7dvdmf4zk7mBS4j4VlkUAN8/2LA4ucYGYe3Kfizeei7VTHkLd2/R9OmYF7Tn+A+PZ
Gyk9h4XNGxfTKFB5U6/ICddnDo57Z1LbcjREKO3Hw/wp5zwTwhbetNG6pJnKQgK9AjfX0zLnE2QQ
jv0x6Nl8roPbkgCe1nbsunvTCikSd/Wvc41dg6M9EVgGX2rHlLb6YBQabH5rynxHHZCXS+4U0dcd
DxIhy94qfa3ovbhpuEBj28VM6HwzyGDoz21HatHXmI8GC3jc8n1ljHp0K1oddu9E8ynj8QA+VZ3x
v5ieBVJbkS5AwImaS3QFAv6MndMFhipzDuBqKXRuyXQTPSzgph18zcixhop2AniuerssYNq6nAsE
nrHtqwJNKrKjGqZeYBYc86D4dlWDs+WrCynGMIXMYO2LnCc6ZPXmHlko+n8y/M3rZEkJu8ikEjcS
VnHzAtVh11XvFUnM+foisk2C0LjFphH3NTXjvahRYKxSnjX9LiV4w6jxdZ5kca6DPnhN7NHaNnnk
sW5yaMJZgm52OL5MOXAHtLc2uLlCjaKts3ehT2IV7TrFT41A3K+h0ijyuYsXn7EuYcF3z9ihAjFT
kYb2E6hKus2zpmkY2PPF2/H7/PxmniatBI0ZC2Q4DNkBkZNxJm7PZkLi0nqVJVAybAmDliP3oaxe
Xgk4FWInCp3IS9QkBpqe9kuNEpj7dS19w6Y9W+ML8iLoO+rJvVGGe0astP0rGR+0G6wcQXZ6J4+n
3kzLszkx6aGjbQ6jWzMPCW1XIaeKoUuYFRazpxwS8vlUR5YcYyTqiGtcwcGHC2Vz3eznyqrbxwxp
dSNw/d5/PrMQy/DL1xg8t3i4Ke5oaJuspEmAFkWJDiN2xpZyfpEVviG3zXfrr6p+YR0kn4r9o3m0
HMjLD2KON8WU0OZHtI3m1obRZQSrpM8kG/72Q3KhrMD0ENtPRMQ+kF9D4mQQ/q1taai42SbyvrJA
4WKeFY57+sUiuUxCloRjPViFlQFrnKMerSn3GeKmhsnxT+sZRRL/CHt5mjbNjxzguu2htli8bvBm
CNPUYGqpuIbuSSan7htmJfAhLXm2kBI2gX7qh+wE7+9O5ImmBjN5U33DjArbBKMXFJVTBjKtrbtX
gMGJlzEu+ghw0j6tRnxr2vtUSzKNhQe3XOuvCmxqGBjbFUlnprMSOyikqA==
`protect end_protected
