--------------------------------------------------------------------------------
-- Engineer:  Luca Caronti    [luca.caronti@studenti.unit.it]
--            Simone Ruffini  [simone.ruffini@tutanota.com]
--
-- Create Date:   05/17/2020 03:21:54 PM
-- Design Name:
-- Module Name:   INT_EMU - Behavioral
-- Project Name:  NORM
--
-- Description: Intermittency emulation core.
-- Details: This entity generates a signal (RST_EMU) used by the test platform
--  as a reset signal. This is generated by comparing a voltage sample to a
--  voltage level selected as the reset threshold.
--
-- Revision:
-- Revision 00 - Luca Caronti
-- * file created
-- Revision 01 - Simone Ruffini
-- * refactoring and generalizatin of the component (input rom is outside of the entity)
-- Additional Comments:
--
--------------------------------------------------------------------------------

----------------------------- PACKAGES/LIBRARIES -------------------------------

library IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.NUMERIC_STD.all;

  -- User libraries
  use work.NORM_PKG.all;

----------------------------- ENTITY -------------------------------------------

entity INT_EMU is
  generic (
    ROMADDR_W           : natural;       -- ROM address bit width
    ROMDOUT_W           : natural;       -- ROM dout bit widht
    NUM_THRESHOLDS      : natural := 1;  -- Number of compared thresholds (the one for RST_EMU is one too)
    SAMPLES_PRESCALER   : natural := 1   -- Sampling from ROM prescaler value (NOTE: > 0)
  );
  port (
    CLK                 : in    std_logic;                                     -- Clock signal
    RST                 : in    std_logic;                                     -- Positive reset
    EN                  : in    std_logic;                                     -- Enable core
    INIT                : in    std_logic;                                     -- Init core
    RST_EMU             : out   std_logic;                                     -- Emulated positive reset
    THRESH_STAT         : out   std_logic_vector(NUM_THRESHOLDS - 1 downto 0); -- Thresholds statuses
    THRESH_VALUES       : in    thresh_values_t(NUM_THRESHOLDS - 1 downto 0);  -- Thresholds values
    RST_EMU_THRESH_INDX : in    natural range 0 to NUM_THRESHOLDS - 1;         -- Index of threshold used for RST_EMU
    ROM_START_ADDR      : in    std_logic_vector(ROMADDR_W - 1 downto 0);      -- ROM start address for sampling
    ROM_OFFSET          : in    natural range 0 to (2 ** ROMADDR_W - 1);       -- ROM last sample, offset from ROM_START_ADDR
    ROM_ADDR            : out   std_logic_vector(ROMADDR_W - 1 downto 0);      -- ROM address
    ROM_DOUT            : in    std_logic_vector(ROMDOUT_W - 1 downto 0)       -- ROM dout
  );
end entity INT_EMU;

----------------------------- ARCHITECTURE -------------------------------------

architecture BEHAVIORAL of INT_EMU is

  --########################### CONSTANTS 1 ####################################

  --########################### TYPES ##########################################

  --########################### FUNCTIONS ######################################

  --########################### CONSTANTS 2 ####################################

  --########################### SIGNALS ########################################

  signal rom_start_addr_samp  : std_logic_vector(ROMADDR_W - 1 downto 0);
  signal rom_offset_samp      : natural range 0 to (2 ** ROMADDR_W - 1);
  signal rom_addr_s           : std_logic_vector(ROMADDR_W - 1 downto 0);
  signal output_comparator    : std_logic_vector(NUM_THRESHOLDS - 1 downto 0);
  signal prescaler_cnt_tc     : std_logic;
  signal prescaler_cnt_init   : std_logic;

  --########################### ARCHITECTURE BEGIN #############################

begin

  assert (SAMPLES_PRESCSLER > 0)
    report "The prescaler for the sampling time must be greater then 0"
    severity failure;

  --########################### ENTITY DEFINITION ##############################

  U_PRESCALER : entity work.cnt
    generic map (
      MAX         => SAMPLES_PRESCALER - 1,
      INIT_VALUE  => SAMPLES_PRESCALER - 1,
      INCREASE_BY => 1
    )
    port map (
      CLK   => CLK,
      RST   => RST,
      INIT  => prescaler_cnt_init,
      CE    => '1',
      TC    => prescaler_cnt_tc,
      VALUE => open
    );

  --########################## OUTPUT PORTS WIRING #############################

  G_COMPARATOR : for i in NUM_THRESHOLDS - 1  downto 0 generate
    output_comparator(i) <= '0' when unsigned(ROM_DOUT) > THRESH_VALUES(i) else
                            '1';
  end generate G_COMPARATOR;

  RESET_EMULATOR <= output_comparator(RST_EMU_THRESH_INDX);

  THRESH_STAT <= output_comparator;

  ROM_ADDR <= rom_addr_s;

  --########################## PROCESSES #######################################

  -- Keep init signal after rst is down for the rest of the clock cycle
  -- this lets PRESCALER_CNT more init time
  P_KEEP_INIT : process (CLK) is
  begin

    if (CLK'event and CLK = '1') then
      prescaler_cnt_init <= '0';
      if (RST = '1') then
        prescaler_cnt_init <= '1';
      end if;
    end if;

  end process P_KEEP_INIT;

  -- Samples rom start address and rom offset
  -- These signals can change only after an init
  P_SAMP : process (CLK, RST) is
  begin

    if (RST = '1') then
      rom_start_addr_samp <= (others => '0');
      rom_offset_samp     <= (others => '0');
    elsif (CLK'event and CLK = '1') then
      if (INIT = '1') then
        rom_start_addr_samp <= ROM_START_ADDR;
        rom_offset_samp     <= ROM_OFFSET;
      end if;
    end if;

  end process P_SAMP;

  -- Calculate rom address, and on overflow start from beginning
  P_ROM_ADDR : process (CLK, RST) is
  begin

    if (RST = '1') then
      rom_s <= (others => '0');
    elsif (CLK'event and CLK = '1') then
      if (INIT = '1') then
        rom_s <= ROM_START_ADDR;
      end if;

      if (EN = '1' AND prescaler_cnt_tc = '1') then
        if (rom_s = std_logic_vector(unsigned(rom_start_addr_samp) + rom_offset_samp)) then
          roms_s <= rom_start_addr_samp;
        else
          rom_s <= std_logic(unsigned(rom_s) + 1);
        end if;
      end if;
    end if;

  end process P_ROM_ADDR;

end architecture BEHAVIORAL;

--------------------------------------------------------------------------------
